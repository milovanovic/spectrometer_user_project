// SPDX-License-Identifier: Apache-2.0

module AXI4HyperSpace(
  input         clock,
  input         reset,
  output        ioMem_0_aw_ready,
  input         ioMem_0_aw_valid,
  input         ioMem_0_aw_bits_id,
  input  [31:0] ioMem_0_aw_bits_addr,
  input  [7:0]  ioMem_0_aw_bits_len,
  input  [2:0]  ioMem_0_aw_bits_size,
  input  [1:0]  ioMem_0_aw_bits_burst,
  input         ioMem_0_aw_bits_lock,
  input  [3:0]  ioMem_0_aw_bits_cache,
  input  [2:0]  ioMem_0_aw_bits_prot,
  input  [3:0]  ioMem_0_aw_bits_qos,
  output        ioMem_0_w_ready,
  input         ioMem_0_w_valid,
  input  [31:0] ioMem_0_w_bits_data,
  input  [3:0]  ioMem_0_w_bits_strb,
  input         ioMem_0_w_bits_last,
  input         ioMem_0_b_ready,
  output        ioMem_0_b_valid,
  output        ioMem_0_b_bits_id,
  output [1:0]  ioMem_0_b_bits_resp,
  output        ioMem_0_ar_ready,
  input         ioMem_0_ar_valid,
  input         ioMem_0_ar_bits_id,
  input  [31:0] ioMem_0_ar_bits_addr,
  input  [7:0]  ioMem_0_ar_bits_len,
  input  [2:0]  ioMem_0_ar_bits_size,
  input  [1:0]  ioMem_0_ar_bits_burst,
  input         ioMem_0_ar_bits_lock,
  input  [3:0]  ioMem_0_ar_bits_cache,
  input  [2:0]  ioMem_0_ar_bits_prot,
  input  [3:0]  ioMem_0_ar_bits_qos,
  input         ioMem_0_r_ready,
  output        ioMem_0_r_valid,
  output        ioMem_0_r_bits_id,
  output [31:0] ioMem_0_r_bits_data,
  output [1:0]  ioMem_0_r_bits_resp,
  output        ioMem_0_r_bits_last,
  output        in_0_ready,
  input         in_0_valid,
  input  [7:0]  in_0_bits_data,
  input         in_0_bits_last,
  input         out_0_ready,
  output        out_0_valid,
  output [15:0] out_0_bits_data,
  output        out_0_bits_last,

  output  [7:0] sram_R0_addr,
  output        sram_R0_clk,
  output        sram_R0_en,
  input  [31:0] sram_R0_data,
  output  [7:0] sram_W0_addr,
  output        sram_W0_en,
  output        sram_W0_clk,
  output [31:0] sram_W0_data
);
  wire  widthAdapter_clock;
  wire  widthAdapter_reset;
  wire  widthAdapter_auto_in_ready;
  wire  widthAdapter_auto_in_valid;
  wire [7:0] widthAdapter_auto_in_bits_data;
  wire  widthAdapter_auto_in_bits_last;
  wire  widthAdapter_auto_out_ready;
  wire  widthAdapter_auto_out_valid;
  wire [31:0] widthAdapter_auto_out_bits_data;
  wire  widthAdapter_auto_out_bits_last;
  reg [7:0] widthAdapter__T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg [7:0] widthAdapter__T_1; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_1;
  reg [7:0] widthAdapter__T_2; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg [1:0] widthAdapter__T_3; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire  widthAdapter__T_4; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire  widthAdapter__T_5; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] widthAdapter__T_6; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] widthAdapter__T_7; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] widthAdapter__GEN_0; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  widthAdapter__T_9; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  widthAdapter__T_10; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  widthAdapter__T_12; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  widthAdapter__T_13; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  widthAdapter__T_15; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  widthAdapter__T_16; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [23:0] widthAdapter__T_18; // @[Cat.scala 29:58]
  wire  widthAdapter_ov0; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  widthAdapter__T_20; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_4;
  reg  widthAdapter__T_21; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_5;
  reg  widthAdapter__T_22; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_6;
  reg [1:0] widthAdapter__T_23; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_7;
  wire  widthAdapter__T_25; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] widthAdapter__T_26; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] widthAdapter__T_27; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] widthAdapter__GEN_4; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  widthAdapter__T_29; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  widthAdapter__T_30; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  widthAdapter__T_32; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  widthAdapter__T_33; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  widthAdapter__T_35; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  widthAdapter__T_36; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [3:0] widthAdapter__T_39; // @[Cat.scala 29:58]
  wire  widthAdapter_ov1; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] widthAdapter__T_44; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_8;
  wire  widthAdapter__T_46; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] widthAdapter__T_47; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] widthAdapter__T_48; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] widthAdapter__GEN_8; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  widthAdapter_ov2; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] widthAdapter__T_64; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_9;
  wire  widthAdapter__T_66; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] widthAdapter__T_67; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] widthAdapter__T_68; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] widthAdapter__GEN_12; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  widthAdapter_ov3; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] widthAdapter__T_84; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_10;
  wire  widthAdapter__T_86; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] widthAdapter__T_87; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] widthAdapter__T_88; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] widthAdapter__GEN_16; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  widthAdapter_ov4; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  widthAdapter__T_101; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  widthAdapter__T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  widthAdapter__T_104; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  widthAdapter__T_105; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  widthAdapter__T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  widthAdapter__T_108; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  widthAdapter__T_109; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  widthAdapter__T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  widthAdapter__T_112; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  widthAdapter__T_113; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  widthAdapter__T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  widthAdapter__T_116; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  fft_clock;
  wire  fft_reset;
  wire  fft_auto_mem_in_aw_ready;
  wire  fft_auto_mem_in_aw_valid;
  wire  fft_auto_mem_in_aw_bits_id;
  wire [29:0] fft_auto_mem_in_aw_bits_addr;
  wire  fft_auto_mem_in_w_ready;
  wire  fft_auto_mem_in_w_valid;
  wire  fft_auto_mem_in_b_ready;
  wire  fft_auto_mem_in_b_valid;
  wire  fft_auto_mem_in_b_bits_id;
  wire  fft_auto_mem_in_ar_ready;
  wire  fft_auto_mem_in_ar_valid;
  wire  fft_auto_mem_in_ar_bits_id;
  wire [29:0] fft_auto_mem_in_ar_bits_addr;
  wire  fft_auto_mem_in_r_ready;
  wire  fft_auto_mem_in_r_valid;
  wire  fft_auto_mem_in_r_bits_id;
  wire [31:0] fft_auto_mem_in_r_bits_data;
  wire  fft_auto_stream_in_ready;
  wire  fft_auto_stream_in_valid;
  wire [31:0] fft_auto_stream_in_bits_data;
  wire  fft_auto_stream_in_bits_last;
  wire  fft_auto_stream_out_ready;
  wire  fft_auto_stream_out_valid;
  wire [31:0] fft_auto_stream_out_bits_data;
  wire  fft_auto_stream_out_bits_last;
  wire  fft_fft_clock;
  wire  fft_fft_reset;
  wire  fft_fft_io_in_ready;
  wire  fft_fft_io_in_valid;
  wire [15:0] fft_fft_io_in_bits_real;
  wire [15:0] fft_fft_io_in_bits_imag;
  wire  fft_fft_io_out_ready;
  wire  fft_fft_io_out_valid;
  wire [15:0] fft_fft_io_out_bits_real;
  wire [15:0] fft_fft_io_out_bits_imag;
  wire  fft_fft_io_lastOut;
  wire  fft_fft_io_lastIn;
  wire  fft_fft_io_busy;
  wire  fft_fft_SDFChainRadix22_clock;
  wire  fft_fft_SDFChainRadix22_reset;
  wire  fft_fft_SDFChainRadix22_io_in_ready;
  wire  fft_fft_SDFChainRadix22_io_in_valid;
  wire [15:0] fft_fft_SDFChainRadix22_io_in_bits_real;
  wire [15:0] fft_fft_SDFChainRadix22_io_in_bits_imag;
  wire  fft_fft_SDFChainRadix22_io_out_ready;
  wire  fft_fft_SDFChainRadix22_io_out_valid;
  wire [15:0] fft_fft_SDFChainRadix22_io_out_bits_real;
  wire [15:0] fft_fft_SDFChainRadix22_io_out_bits_imag;
  wire  fft_fft_SDFChainRadix22_io_lastOut;
  wire  fft_fft_SDFChainRadix22_io_lastIn;
  wire  fft_fft_SDFChainRadix22_io_busy;
  wire  fft_fft_SDFChainRadix22_sdf_stages_0_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_0_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_0_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_0_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_47; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_49; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_52; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_54; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_56; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_59; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_30; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_32; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_35; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_37; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_39; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_0__T_42; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_0_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_1_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_1_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_1_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_1_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_50; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_52; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_55; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_57; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_59; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_62; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_33; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_35; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_38; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_40; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_42; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_1__T_45; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_1_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_2_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_2_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_2_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_2_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_56; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_58; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_61; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_63; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_65; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_68; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_39; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_41; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_44; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_46; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_48; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_2__T_51; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_2_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_3_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_3_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_3_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_3_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_68; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_70; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_73; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_75; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_77; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_80; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_51; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_53; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_56; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_58; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_60; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_3__T_63; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_3_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_4_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_4_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_4_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_4_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_92; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_94; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_97; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_99; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_101; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_104; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_75; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_77; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_80; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_82; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_84; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_4__T_87; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_4_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_5_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_5_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_5_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_5_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_140; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_142; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_145; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_147; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_149; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_152; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_123; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_125; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_128; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_130; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_132; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_5__T_135; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_5_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_6_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_6_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_6_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_6_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_236; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_238; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_241; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_243; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_245; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_248; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_114_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_114_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_117_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_117_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_120_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_120_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_123_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_123_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_126_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_126_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_129_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_129_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_132_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_132_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_135_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_135_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_138_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_138_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_141_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_141_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_144_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_144_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_147_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_147_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_150_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_150_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_153_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_153_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_156_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_156_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_159_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_159_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_162_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_162_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_165_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_165_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_168_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_168_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_171_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_171_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_174_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_174_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_177_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_177_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_180_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_180_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_183_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_183_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_186_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_186_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_189_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_189_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_192_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_192_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_195_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_195_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_198_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_198_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_201_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_201_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_204_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_204_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_207_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_207_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_219; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_221; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_224; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_226; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_228; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_6__T_231; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_6_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_7_clock;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_7_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_7_io_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_7_load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_428; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_430; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_433; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_435; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_437; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_440; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_114_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_114_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_117_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_117_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_120_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_120_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_123_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_123_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_126_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_126_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_129_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_129_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_132_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_132_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_135_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_135_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_138_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_138_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_141_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_141_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_144_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_144_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_147_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_147_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_150_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_150_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_153_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_153_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_156_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_156_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_159_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_159_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_162_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_162_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_165_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_165_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_168_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_168_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_171_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_171_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_174_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_174_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_177_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_177_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_180_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_180_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_183_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_183_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_186_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_186_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_189_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_189_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_192_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_192_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_195_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_195_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_198_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_198_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_201_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_201_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_204_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_204_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_207_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_207_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_210_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_210_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_213_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_213_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_216_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_216_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_219_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_219_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_222_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_222_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_225_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_225_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_228_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_228_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_231_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_231_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_234_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_234_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_237_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_237_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_240_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_240_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_243_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_243_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_246_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_246_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_249_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_249_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_252_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_252_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_255_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_255_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_258_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_258_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_261_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_261_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_264_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_264_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_267_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_267_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_270_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_270_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_273_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_273_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_276_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_276_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_279_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_279_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_282_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_282_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_285_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_285_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_288_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_288_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_291_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_291_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_294_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_294_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_297_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_297_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_300_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_300_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_303_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_303_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_306_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_306_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_309_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_309_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_312_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_312_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_315_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_315_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_318_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_318_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_321_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_321_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_324_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_324_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_327_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_327_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_330_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_330_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_333_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_333_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_336_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_336_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_339_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_339_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_342_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_342_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_345_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_345_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_348_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_348_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_351_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_351_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_354_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_354_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_357_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_357_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_360_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_360_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_363_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_363_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_366_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_366_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_369_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_369_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_372_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_372_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_375_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_375_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_378_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_378_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_381_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_381_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_384_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_384_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_387_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_387_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_390_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_513;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_390_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_514;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_393_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_515;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_393_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_516;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_396_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_517;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_396_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_518;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_399_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_519;
  reg [15:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_399_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_520;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_411; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_413; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_416; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_418; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_420; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_7__T_423; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_7_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_clock;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_reset;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_io_in_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_io_in_imag;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_io_out_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_io_out_imag;
  wire [8:0] fft_fft_SDFChainRadix22_sdf_stages_8_io_cntr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_io_en;
  wire [7:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_addr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_clk;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_data_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_data_imag;
  wire [7:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_addr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_clk;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_data_real;
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_data_imag;
  wire [7:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_addr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_clk;
  wire [31:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_data;
  wire [7:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_addr;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_en;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_clk;
  wire [31:0] fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_data;
  wire  fft_fft_SDFChainRadix22_sdf_stages_8_load_input; // @[UIntTypeClass.scala 52:47]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_feedback_real; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_57; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_59; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_62; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_feedback_imag; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_64; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_66; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_69; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [7:0] fft_fft_SDFChainRadix22_sdf_stages_8_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_521;
  wire [7:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_22; // @[Counter.scala 39:22]
  reg [7:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_26; // @[Reg.scala 27:20]
  reg [31:0] _RAND_522;
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_40; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_42; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_45; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_47; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_49; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] fft_fft_SDFChainRadix22_sdf_stages_8__T_52; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] fft_fft_SDFChainRadix22_sdf_stages_8_butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [1:0] fft_fft_SDFChainRadix22_state; // @[SDFChainRadix22.scala 56:22]
  reg [31:0] _RAND_523;
  reg  fft_fft_SDFChainRadix22_initialOutDone; // @[SDFChainRadix22.scala 59:31]
  reg [31:0] _RAND_524;
  reg [9:0] fft_fft_SDFChainRadix22_cnt; // @[SDFChainRadix22.scala 60:20]
  reg [31:0] _RAND_525;
  wire  fft_fft_SDFChainRadix22__T_46; // @[Decoupled.scala 40:37]
  wire  fft_fft_SDFChainRadix22_fireLast; // @[SDFChainRadix22.scala 79:28]
  wire [8:0] fft_fft_SDFChainRadix22__T_48; // @[SDFChainRadix22.scala 81:45]
  wire [3:0] fft_fft_SDFChainRadix22__T_49;
  wire  fft_fft_SDFChainRadix22__T_53; // @[Conditional.scala 37:30]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_0; // @[SDFChainRadix22.scala 90:27]
  wire  fft_fft_SDFChainRadix22__T_56; // @[Conditional.scala 37:30]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_1; // @[SDFChainRadix22.scala 93:23]
  wire  fft_fft_SDFChainRadix22__T_57; // @[Conditional.scala 37:30]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_2; // @[SDFChainRadix22.scala 98:25]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_3; // @[Conditional.scala 39:67]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_4; // @[Conditional.scala 39:67]
  wire [1:0] fft_fft_SDFChainRadix22_state_next; // @[Conditional.scala 40:58]
  reg [8:0] fft_fft_SDFChainRadix22_cntValidOut; // @[SDFChainRadix22.scala 106:28]
  reg [31:0] _RAND_526;
  wire [9:0] fft_fft_SDFChainRadix22__T_59; // @[SDFChainRadix22.scala 111:44]
  wire [9:0] fft_fft_SDFChainRadix22__GEN_2109; // @[SDFChainRadix22.scala 111:29]
  wire  fft_fft_SDFChainRadix22__T_60; // @[SDFChainRadix22.scala 111:29]
  wire  fft_fft_SDFChainRadix22__T_61; // @[Decoupled.scala 40:37]
  wire  fft_fft_SDFChainRadix22_pktEnd; // @[SDFChainRadix22.scala 111:52]
  wire  fft_fft_SDFChainRadix22__T_62; // @[SDFChainRadix22.scala 114:20]
  wire [8:0] fft_fft_SDFChainRadix22_cntr_wires_0; // @[SDFChainRadix22.scala 52:24 SDFChainRadix22.scala 185:29]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_20; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_21; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_22; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_23; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_24; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_25; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_26; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] fft_fft_SDFChainRadix22__GEN_27; // @[SDFChainRadix22.scala 126:79]
  wire [9:0] fft_fft_SDFChainRadix22__GEN_2110; // @[SDFChainRadix22.scala 126:79]
  wire  fft_fft_SDFChainRadix22__T_76; // @[SDFChainRadix22.scala 130:31]
  wire  fft_fft_SDFChainRadix22__T_77; // @[SDFChainRadix22.scala 130:42]
  wire [8:0] fft_fft_SDFChainRadix22__T_80; // @[SDFChainRadix22.scala 134:32]
  wire  fft_fft_SDFChainRadix22__T_83; // @[SDFChainRadix22.scala 144:90]
  wire  fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 173:54]
  wire  fft_fft_SDFChainRadix22_enableInit; // @[SDFChainRadix22.scala 173:33]
  wire [9:0] fft_fft_SDFChainRadix22__T_125; // @[SDFChainRadix22.scala 179:16]
  wire [9:0] fft_fft_SDFChainRadix22__T_145; // @[SDFChainRadix22.scala 193:37]
  wire  fft_fft_SDFChainRadix22__T_146; // @[SDFChainRadix22.scala 193:22]
  wire  fft_fft_SDFChainRadix22__T_147; // @[SDFChainRadix22.scala 193:44]
  wire  fft_fft_SDFChainRadix22__GEN_45; // @[SDFChainRadix22.scala 196:36]
  wire  fft_fft_SDFChainRadix22__GEN_46; // @[SDFChainRadix22.scala 193:60]
  wire [8:0] fft_fft_SDFChainRadix22__T_166; // @[SDFChainRadix22.scala 224:38]
  wire  fft_fft_SDFChainRadix22__T_167; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_171; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] fft_fft_SDFChainRadix22__T_173; // @[SDFChainRadix22.scala 224:38]
  wire [1:0] fft_fft_SDFChainRadix22__T_174; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_178; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] fft_fft_SDFChainRadix22__T_180; // @[SDFChainRadix22.scala 224:38]
  wire [2:0] fft_fft_SDFChainRadix22__T_181; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_185; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] fft_fft_SDFChainRadix22__T_187; // @[SDFChainRadix22.scala 224:38]
  wire [3:0] fft_fft_SDFChainRadix22__T_188; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_192; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] fft_fft_SDFChainRadix22__T_194; // @[SDFChainRadix22.scala 224:38]
  wire [4:0] fft_fft_SDFChainRadix22__T_195; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_199; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] fft_fft_SDFChainRadix22__T_201; // @[SDFChainRadix22.scala 224:38]
  wire [5:0] fft_fft_SDFChainRadix22__T_202; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_206; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] fft_fft_SDFChainRadix22__T_208; // @[SDFChainRadix22.scala 224:38]
  wire [6:0] fft_fft_SDFChainRadix22__T_209; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_213; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] fft_fft_SDFChainRadix22__T_215; // @[SDFChainRadix22.scala 224:38]
  wire [7:0] fft_fft_SDFChainRadix22__T_216; // @[SDFChainRadix22.scala 224:92]
  wire [8:0] fft_fft_SDFChainRadix22__T_220; // @[SDFChainRadix22.scala 224:68]
  wire [2:0] fft_fft_SDFChainRadix22__T_255;
  wire [1:0] fft_fft_SDFChainRadix22__GEN_52; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_53; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_54; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_55; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] fft_fft_SDFChainRadix22__GEN_56; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_59; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_60; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_61; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_62; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_63; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22_twiddles_1_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] fft_fft_SDFChainRadix22__T_261; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_0_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_0_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  wire [16:0] fft_fft_SDFChainRadix22__T_262; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22__T_263; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2112; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_264; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2113; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_265; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2114; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_266; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] fft_fft_SDFChainRadix22__T_267; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_268; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_274; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_275; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] fft_fft_SDFChainRadix22__T_278; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_279; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22__T_286; // @[SDFChainRadix22.scala 328:32]
  wire  fft_fft_SDFChainRadix22__T_287; // @[SDFChainRadix22.scala 328:78]
  wire  fft_fft_SDFChainRadix22__T_288; // @[SDFChainRadix22.scala 328:65]
  wire  fft_fft_SDFChainRadix22__T_289; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_1_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] fft_fft_SDFChainRadix22__T_295; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_1_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [4:0] fft_fft_SDFChainRadix22__T_387;
  wire [3:0] fft_fft_SDFChainRadix22__GEN_82; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_83; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_84; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_85; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_86; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_87; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_88; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_89; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_90; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_91; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_92; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_93; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_94; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_95; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_96; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_97; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_98; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_99; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_100; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_101; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_102; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_103; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] fft_fft_SDFChainRadix22__GEN_104; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_107; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_108; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_109; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_110; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_111; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_112; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_113; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_114; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_115; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_116; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_117; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_118; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_119; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_120; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_121; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_122; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_123; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_124; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_125; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_126; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_127; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_128; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_129; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_130; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_131; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_132; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_133; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_134; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_135; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22_twiddles_3_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] fft_fft_SDFChainRadix22__T_393; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_2_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_2_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [16:0] fft_fft_SDFChainRadix22__T_394; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22__T_395; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2115; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_396; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2116; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_397; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2117; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_398; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] fft_fft_SDFChainRadix22__T_399; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_400; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_406; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_407; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] fft_fft_SDFChainRadix22__T_410; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_411; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22__T_418; // @[SDFChainRadix22.scala 328:32]
  wire  fft_fft_SDFChainRadix22__T_419; // @[SDFChainRadix22.scala 328:78]
  wire  fft_fft_SDFChainRadix22__T_420; // @[SDFChainRadix22.scala 328:65]
  wire  fft_fft_SDFChainRadix22__T_421; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_3_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] fft_fft_SDFChainRadix22__T_427; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_3_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [6:0] fft_fft_SDFChainRadix22__T_759;
  wire [5:0] fft_fft_SDFChainRadix22__GEN_202; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_203; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_204; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_205; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_206; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_207; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_208; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_209; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_210; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_211; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_212; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_213; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_214; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_215; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_216; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_217; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_218; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_219; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_220; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_221; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_222; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_223; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_224; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_225; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_226; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_227; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_228; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_229; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_230; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_231; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_232; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_233; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_234; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_235; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_236; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_237; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_238; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_239; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_240; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_241; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_242; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_243; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_244; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_245; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_246; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_247; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_248; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_249; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_250; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_251; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_252; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_253; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_254; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_255; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_256; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_257; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_258; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_259; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_260; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_261; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_262; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_263; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_264; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_265; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_266; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_267; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_268; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_269; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_270; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_271; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_272; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_273; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_274; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_275; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_276; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_277; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_278; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_279; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_280; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_281; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_282; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_283; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_284; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_285; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_286; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_287; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_288; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_289; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_290; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_291; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_292; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_293; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_294; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_295; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] fft_fft_SDFChainRadix22__GEN_296; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_299; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_300; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_301; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_302; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_303; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_304; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_305; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_306; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_307; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_308; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_309; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_310; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_311; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_312; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_313; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_314; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_315; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_316; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_317; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_318; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_319; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_320; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_321; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_322; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_323; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_324; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_325; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_326; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_327; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_328; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_329; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_330; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_331; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_332; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_333; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_334; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_335; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_336; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_337; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_338; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_339; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_340; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_341; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_342; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_343; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_344; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_345; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_346; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_347; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_348; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_349; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_350; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_351; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_352; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_353; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_354; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_355; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_356; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_357; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_358; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_359; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_360; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_361; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_362; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_363; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_364; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_365; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_366; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_367; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_368; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_369; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_370; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_371; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_372; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_373; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_374; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_375; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_376; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_377; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_378; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_379; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_380; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_381; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_382; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_383; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_384; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_385; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_386; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_387; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_388; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_389; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_390; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_391; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_392; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_393; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_394; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_395; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_396; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_397; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_398; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_399; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_400; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_401; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_402; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_403; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_404; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_405; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_406; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_407; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_408; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_409; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_410; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_411; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_412; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_413; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_414; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_415; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_416; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_417; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_418; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_419; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_420; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_421; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_422; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_423; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22_twiddles_5_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] fft_fft_SDFChainRadix22__T_765; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_4_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_4_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [16:0] fft_fft_SDFChainRadix22__T_766; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22__T_767; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2118; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_768; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2119; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_769; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2120; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_770; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] fft_fft_SDFChainRadix22__T_771; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_772; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_778; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_779; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] fft_fft_SDFChainRadix22__T_782; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_783; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22__T_790; // @[SDFChainRadix22.scala 328:32]
  wire  fft_fft_SDFChainRadix22__T_791; // @[SDFChainRadix22.scala 328:78]
  wire  fft_fft_SDFChainRadix22__T_792; // @[SDFChainRadix22.scala 328:65]
  wire  fft_fft_SDFChainRadix22__T_793; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_5_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] fft_fft_SDFChainRadix22__T_799; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_5_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_682; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_683; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_684; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_685; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_686; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_687; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_688; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_689; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_690; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_691; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_692; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_693; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_694; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_695; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_696; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_697; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_698; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_699; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_700; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_701; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_702; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_703; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_704; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_705; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_706; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_707; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_708; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_709; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_710; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_711; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_712; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_713; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_714; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_715; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_716; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_717; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_718; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_719; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_720; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_721; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_722; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_723; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_724; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_725; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_726; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_727; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_728; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_729; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_730; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_731; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_732; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_733; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_734; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_735; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_736; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_737; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_738; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_739; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_740; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_741; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_742; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_743; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_744; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_745; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_746; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_747; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_748; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_749; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_750; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_751; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_752; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_753; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_754; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_755; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_756; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_757; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_758; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_759; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_760; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_761; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_762; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_763; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_764; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_765; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_766; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_767; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_768; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_769; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_770; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_771; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_772; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_773; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_774; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_775; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_776; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_777; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_778; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_779; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_780; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_781; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_782; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_783; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_784; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_785; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_786; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_787; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_788; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_789; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_790; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_791; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_792; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_793; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_794; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_795; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_796; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_797; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_798; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_799; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_800; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_801; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_802; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_803; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_804; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_805; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_806; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_807; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_808; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_809; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_810; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_811; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_812; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_813; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_814; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_815; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_816; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_817; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_818; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_819; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_820; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_821; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_822; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_823; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_824; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_825; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_826; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_827; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_828; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_829; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_830; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_831; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_832; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_833; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_834; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_835; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_836; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_837; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_838; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_839; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_840; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_841; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_842; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_843; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_844; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_845; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_846; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_847; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_848; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_849; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_850; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_851; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_852; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_853; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_854; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_855; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_856; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_857; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_858; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_859; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_860; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_861; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_862; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_863; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_864; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_865; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_866; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_867; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_868; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_869; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_870; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_871; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_872; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_873; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_874; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_875; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_876; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_877; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_878; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_879; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_880; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_881; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_882; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_883; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_884; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_885; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_886; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_887; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_888; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_889; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_890; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_891; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_892; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_893; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_894; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_895; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_896; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_897; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_898; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_899; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_900; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_901; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_902; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_903; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_904; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_905; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_906; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_907; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_908; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_909; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_910; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_911; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_912; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_913; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_914; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_915; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_916; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_917; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_918; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_919; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_920; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_921; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_922; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_923; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_924; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_925; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_926; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_927; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_928; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_929; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_930; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_931; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_932; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_933; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_934; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_935; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_936; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_937; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_938; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_939; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_940; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_941; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_942; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_943; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_944; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_945; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_946; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_947; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_948; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_949; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_950; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_951; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_952; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_953; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_954; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_955; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_956; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_957; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_958; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_959; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_960; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_961; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_962; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_963; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_964; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_965; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_966; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_967; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_968; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_969; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_970; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_971; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_972; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_973; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_974; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_975; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_976; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_977; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_978; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_979; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_980; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_981; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_982; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_983; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_984; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_985; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_986; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_987; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_988; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_989; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_990; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_991; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_992; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_993; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_994; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_995; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_996; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_997; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_998; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_999; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1000; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1001; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1002; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1003; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1004; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1005; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1006; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1007; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1008; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1009; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1010; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1011; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1012; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1013; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1014; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1015; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1016; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1017; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1018; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1019; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1020; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1021; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1022; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1023; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1024; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1025; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1026; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1027; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1028; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1029; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1030; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1031; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1032; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1033; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1034; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1035; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1036; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1037; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1038; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1039; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1040; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1041; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1042; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1043; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1044; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1045; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1046; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1047; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1048; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1049; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1050; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1051; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1052; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1053; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1054; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1055; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1056; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1057; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1058; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1059; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1060; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1061; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1062; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1063; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] fft_fft_SDFChainRadix22__GEN_1064; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1067; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1068; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1069; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1070; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1071; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1072; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1073; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1074; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1075; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1076; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1077; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1078; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1079; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1080; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1081; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1082; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1083; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1084; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1085; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1086; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1087; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1088; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1089; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1090; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1091; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1092; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1093; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1094; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1095; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1096; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1097; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1098; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1099; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1100; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1101; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1102; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1103; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1104; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1105; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1106; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1107; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1108; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1109; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1110; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1111; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1112; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1113; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1114; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1115; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1116; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1117; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1118; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1119; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1120; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1121; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1122; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1123; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1124; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1125; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1126; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1127; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1128; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1129; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1130; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1131; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1132; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1133; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1134; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1135; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1136; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1137; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1138; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1139; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1140; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1141; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1142; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1143; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1144; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1145; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1146; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1147; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1148; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1149; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1150; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1151; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1152; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1153; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1154; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1155; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1156; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1157; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1158; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1159; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1160; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1161; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1162; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1163; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1164; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1165; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1166; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1167; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1168; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1169; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1170; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1171; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1172; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1173; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1174; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1175; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1176; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1177; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1178; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1179; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1180; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1181; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1182; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1183; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1184; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1185; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1186; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1187; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1188; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1189; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1190; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1191; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1192; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1193; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1194; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1195; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1196; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1197; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1198; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1199; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1200; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1201; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1202; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1203; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1204; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1205; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1206; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1207; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1208; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1209; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1210; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1211; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1212; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1213; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1214; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1215; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1216; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1217; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1218; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1219; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1220; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1221; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1222; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1223; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1224; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1225; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1226; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1227; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1228; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1229; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1230; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1231; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1232; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1233; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1234; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1235; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1236; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1237; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1238; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1239; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1240; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1241; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1242; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1243; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1244; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1245; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1246; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1247; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1248; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1249; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1250; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1251; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1252; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1253; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1254; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1255; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1256; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1257; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1258; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1259; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1260; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1261; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1262; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1263; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1264; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1265; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1266; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1267; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1268; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1269; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1270; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1271; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1272; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1273; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1274; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1275; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1276; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1277; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1278; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1279; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1280; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1281; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1282; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1283; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1284; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1285; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1286; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1287; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1288; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1289; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1290; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1291; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1292; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1293; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1294; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1295; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1296; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1297; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1298; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1299; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1300; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1301; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1302; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1303; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1304; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1305; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1306; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1307; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1308; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1309; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1310; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1311; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1312; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1313; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1314; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1315; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1316; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1317; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1318; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1319; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1320; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1321; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1322; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1323; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1324; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1325; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1326; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1327; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1328; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1329; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1330; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1331; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1332; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1333; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1334; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1335; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1336; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1337; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1338; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1339; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1340; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1341; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1342; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1343; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1344; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1345; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1346; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1347; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1348; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1349; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1350; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1351; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1352; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1353; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1354; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1355; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1356; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1357; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1358; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1359; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1360; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1361; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1362; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1363; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1364; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1365; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1366; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1367; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1368; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1369; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1370; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1371; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1372; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1373; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1374; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1375; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1376; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1377; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1378; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1379; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1380; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1381; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1382; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1383; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1384; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1385; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1386; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1387; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1388; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1389; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1390; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1391; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1392; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1393; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1394; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1395; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1396; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1397; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1398; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1399; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1400; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1401; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1402; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1403; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1404; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1405; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1406; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1407; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1408; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1409; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1410; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1411; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1412; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1413; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1414; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1415; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1416; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1417; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1418; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1419; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1420; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1421; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1422; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1423; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1424; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1425; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1426; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1427; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1428; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1429; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1430; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1431; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1432; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1433; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1434; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1435; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1436; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1437; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1438; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1439; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1440; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1441; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1442; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1443; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1444; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1445; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1446; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1447; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1448; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1449; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1450; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1451; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1452; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1453; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1454; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1455; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1456; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1457; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1458; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1459; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1460; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1461; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1462; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1463; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1464; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1465; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1466; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1467; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1468; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1469; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1470; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1471; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1472; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1473; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1474; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1475; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1476; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1477; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1478; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1479; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1480; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1481; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1482; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1483; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1484; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1485; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1486; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1487; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1488; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1489; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1490; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1491; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1492; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1493; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1494; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1495; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1496; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1497; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1498; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1499; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1500; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1501; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1502; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1503; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1504; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1505; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1506; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1507; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1508; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1509; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1510; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1511; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1512; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1513; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1514; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1515; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1516; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1517; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1518; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1519; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1520; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1521; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1522; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1523; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1524; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1525; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1526; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1527; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1528; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1529; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1530; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1531; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1532; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1533; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1534; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1535; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1536; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1537; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1538; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1539; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1540; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1541; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1542; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1543; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1544; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1545; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1546; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1547; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1548; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1549; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1550; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1551; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1552; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1553; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1554; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1555; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1556; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1557; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1558; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1559; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1560; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1561; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1562; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1563; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1564; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1565; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1566; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1567; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1568; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1569; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1570; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1571; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1572; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1573; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1574; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_1575; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] fft_fft_SDFChainRadix22_twiddles_7_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] fft_fft_SDFChainRadix22__T_2096; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_6_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_6_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [16:0] fft_fft_SDFChainRadix22__T_2097; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] fft_fft_SDFChainRadix22__T_2098; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2121; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_2099; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2122; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_2100; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] fft_fft_SDFChainRadix22__GEN_2123; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] fft_fft_SDFChainRadix22__T_2101; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] fft_fft_SDFChainRadix22__T_2102; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_2103; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] fft_fft_SDFChainRadix22__T_2109; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_2110; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] fft_fft_SDFChainRadix22__T_2113; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] fft_fft_SDFChainRadix22__T_2114; // @[FixedPointTypeClass.scala 176:41]
  wire  fft_fft_SDFChainRadix22__T_2121; // @[SDFChainRadix22.scala 328:32]
  wire  fft_fft_SDFChainRadix22__T_2122; // @[SDFChainRadix22.scala 328:78]
  wire  fft_fft_SDFChainRadix22__T_2123; // @[SDFChainRadix22.scala 328:65]
  wire  fft_fft_SDFChainRadix22__T_2124; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_7_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] fft_fft_SDFChainRadix22__T_2130; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_7_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2091; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2092; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2093; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2094; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2095; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2096; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2097; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2098; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2099; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2100; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2101; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2102; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2103; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2104; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_8_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2105; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] fft_fft_SDFChainRadix22_outputWires_8_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] fft_fft_SDFChainRadix22__GEN_2106; // @[SDFChainRadix22.scala 364:24]
  wire  fft_fft_SDFChainRadix22__T_2140; // @[SDFChainRadix22.scala 368:33]
  wire  fft_fft_SDFChainRadix22__T_2141; // @[SDFChainRadix22.scala 368:127]
  wire  fft_fft_SDFChainRadix22__T_2142; // @[SDFChainRadix22.scala 368:117]
  wire [29:0] fft_fft_SDFChainRadix22__GEN_2124; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] fft_fft_SDFChainRadix22__GEN_2107; // @[SDFChainRadix22.scala 375:33]
  wire [29:0] fft_fft_SDFChainRadix22__GEN_2125; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] fft_fft_SDFChainRadix22__GEN_2108; // @[SDFChainRadix22.scala 375:33]
  wire [17:0] fft_fft_SDFChainRadix22__GEN_2126; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 396:27]
  wire [17:0] fft_fft_SDFChainRadix22__GEN_2128; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 397:27]
  wire [31:0] fft_fft__T_152; // @[FixedPointTypeClass.scala 42:59]
  wire [31:0] fft_fft__T_153; // @[FixedPointTypeClass.scala 42:59]
  wire [17:0] fft_fft__GEN_526; // @[SDFFFT.scala 301:31 SDFFFT.scala 309:21]
  wire [17:0] fft_fft__GEN_528; // @[SDFFFT.scala 302:31 SDFFFT.scala 309:21]
  wire  fft_Queue_clock;
  wire  fft_Queue_reset;
  wire  fft_Queue_io_enq_ready;
  wire  fft_Queue_io_enq_valid;
  wire  fft_Queue_io_enq_bits_read;
  wire [31:0] fft_Queue_io_enq_bits_data;
  wire  fft_Queue_io_enq_bits_extra;
  wire  fft_Queue_io_deq_ready;
  wire  fft_Queue_io_deq_valid;
  wire  fft_Queue_io_deq_bits_read;
  wire [31:0] fft_Queue_io_deq_bits_data;
  wire  fft_Queue_io_deq_bits_extra;
  reg  fft_Queue__T_read [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_527;
  wire  fft_Queue__T_read__T_18_data; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_read__T_18_addr; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_read__T_10_data; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_read__T_10_addr; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_read__T_10_mask; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_read__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] fft_Queue__T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_528;
  wire [31:0] fft_Queue__T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] fft_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  fft_Queue__T_extra [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_529;
  wire  fft_Queue__T_extra__T_18_data; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_extra__T_18_addr; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_extra__T_10_data; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_extra__T_10_addr; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_extra__T_10_mask; // @[Decoupled.scala 209:24]
  wire  fft_Queue__T_extra__T_10_en; // @[Decoupled.scala 209:24]
  reg  fft_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_530;
  reg  fft_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_531;
  reg  fft_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_532;
  wire  fft_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  fft_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  fft_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  fft_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  fft_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  fft_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  fft_Queue__T_12; // @[Counter.scala 39:22]
  wire  fft_Queue__T_14; // @[Counter.scala 39:22]
  wire  fft_Queue__T_15; // @[Decoupled.scala 227:16]
  reg  fft_busy; // @[FFTBlock.scala 63:34]
  reg [31:0] _RAND_533;
  wire  fft__T_2; // @[RegisterRouter.scala 40:39]
  wire  fft__T_4; // @[RegisterRouter.scala 42:29]
  wire  fft__T_47_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] fft__T_11; // @[RegisterRouter.scala 48:19]
  wire [27:0] fft__T_45; // @[RegisterRouter.scala 52:27]
  wire [5:0] fft__T_1_bits_index; // @[RegisterRouter.scala 37:18 RegisterRouter.scala 52:19]
  wire  fft__T_53; // @[RegisterRouter.scala 59:16]
  wire  fft__T_5; // @[RegisterRouter.scala 42:26]
  wire  fft__T_171; // @[RegisterRouter.scala 59:16]
  wire  fft__T_172_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  fft__T_172_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  fft__T_175; // @[RegisterRouter.scala 65:29]
  wire  mag_clock;
  wire  mag_reset;
  wire  mag_auto_mem_in_aw_ready;
  wire  mag_auto_mem_in_aw_valid;
  wire  mag_auto_mem_in_aw_bits_id;
  wire [29:0] mag_auto_mem_in_aw_bits_addr;
  wire  mag_auto_mem_in_w_ready;
  wire  mag_auto_mem_in_w_valid;
  wire [31:0] mag_auto_mem_in_w_bits_data;
  wire [3:0] mag_auto_mem_in_w_bits_strb;
  wire  mag_auto_mem_in_b_ready;
  wire  mag_auto_mem_in_b_valid;
  wire  mag_auto_mem_in_b_bits_id;
  wire  mag_auto_mem_in_ar_ready;
  wire  mag_auto_mem_in_ar_valid;
  wire  mag_auto_mem_in_ar_bits_id;
  wire [29:0] mag_auto_mem_in_ar_bits_addr;
  wire [2:0] mag_auto_mem_in_ar_bits_size;
  wire  mag_auto_mem_in_r_ready;
  wire  mag_auto_mem_in_r_valid;
  wire  mag_auto_mem_in_r_bits_id;
  wire [31:0] mag_auto_mem_in_r_bits_data;
  wire  mag_auto_master_out_ready;
  wire  mag_auto_master_out_valid;
  wire [15:0] mag_auto_master_out_bits_data;
  wire  mag_auto_master_out_bits_last;
  wire  mag_auto_slave_in_ready;
  wire  mag_auto_slave_in_valid;
  wire [31:0] mag_auto_slave_in_bits_data;
  wire  mag_auto_slave_in_bits_last;
  wire  mag_logMagMux_clock;
  wire  mag_logMagMux_reset;
  wire  mag_logMagMux_io_in_ready;
  wire  mag_logMagMux_io_in_valid;
  wire [15:0] mag_logMagMux_io_in_bits_real;
  wire [15:0] mag_logMagMux_io_in_bits_imag;
  wire  mag_logMagMux_io_lastIn;
  wire  mag_logMagMux_io_out_ready;
  wire  mag_logMagMux_io_out_valid;
  wire [15:0] mag_logMagMux_io_out_bits;
  wire [1:0] mag_logMagMux_io_sel;
  wire  mag_logMagMux_io_lastOut;
  wire  mag_logMagMux_magModule_clock;
  wire  mag_logMagMux_magModule_reset;
  wire  mag_logMagMux_magModule_io_in_ready;
  wire  mag_logMagMux_magModule_io_in_valid;
  wire [15:0] mag_logMagMux_magModule_io_in_bits_real;
  wire [15:0] mag_logMagMux_magModule_io_in_bits_imag;
  wire  mag_logMagMux_magModule_io_lastIn;
  wire  mag_logMagMux_magModule_io_out_ready;
  wire  mag_logMagMux_magModule_io_out_valid;
  wire [15:0] mag_logMagMux_magModule_io_out_bits;
  wire [1:0] mag_logMagMux_magModule_io_sel;
  wire  mag_logMagMux_magModule_io_lastOut;
  wire  mag_logMagMux_magModule_Queue_clock;
  wire  mag_logMagMux_magModule_Queue_reset;
  wire  mag_logMagMux_magModule_Queue_io_enq_ready;
  wire  mag_logMagMux_magModule_Queue_io_enq_valid;
  wire [15:0] mag_logMagMux_magModule_Queue_io_enq_bits;
  wire  mag_logMagMux_magModule_Queue_io_deq_ready;
  wire  mag_logMagMux_magModule_Queue_io_deq_valid;
  wire [15:0] mag_logMagMux_magModule_Queue_io_deq_bits;
  reg [15:0] mag_logMagMux_magModule_Queue__T [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_534;
  wire [15:0] mag_logMagMux_magModule_Queue__T__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] mag_logMagMux_magModule_Queue__T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] mag_logMagMux_magModule_Queue__T__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] mag_logMagMux_magModule_Queue__T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  mag_logMagMux_magModule_Queue__T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  mag_logMagMux_magModule_Queue__T__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] mag_logMagMux_magModule_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_535;
  reg [1:0] mag_logMagMux_magModule_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_536;
  reg  mag_logMagMux_magModule_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_537;
  wire  mag_logMagMux_magModule_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  mag_logMagMux_magModule_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  mag_logMagMux_magModule_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  mag_logMagMux_magModule_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  mag_logMagMux_magModule_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  mag_logMagMux_magModule_Queue__T_8; // @[Decoupled.scala 40:37]
  wire [1:0] mag_logMagMux_magModule_Queue__T_12; // @[Counter.scala 39:22]
  wire [1:0] mag_logMagMux_magModule_Queue__T_14; // @[Counter.scala 39:22]
  wire  mag_logMagMux_magModule_Queue__T_15; // @[Decoupled.scala 227:16]
  wire  mag_logMagMux_magModule_Queue_1_clock;
  wire  mag_logMagMux_magModule_Queue_1_reset;
  wire  mag_logMagMux_magModule_Queue_1_io_enq_ready;
  wire  mag_logMagMux_magModule_Queue_1_io_enq_valid;
  wire  mag_logMagMux_magModule_Queue_1_io_enq_bits;
  wire  mag_logMagMux_magModule_Queue_1_io_deq_ready;
  wire  mag_logMagMux_magModule_Queue_1_io_deq_valid;
  wire  mag_logMagMux_magModule_Queue_1_io_deq_bits;
  reg  mag_logMagMux_magModule_Queue_1__T [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_538;
  wire  mag_logMagMux_magModule_Queue_1__T__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] mag_logMagMux_magModule_Queue_1__T__T_18_addr; // @[Decoupled.scala 209:24]
  wire  mag_logMagMux_magModule_Queue_1__T__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] mag_logMagMux_magModule_Queue_1__T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  mag_logMagMux_magModule_Queue_1__T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  mag_logMagMux_magModule_Queue_1__T__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] mag_logMagMux_magModule_Queue_1_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_539;
  reg [1:0] mag_logMagMux_magModule_Queue_1_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_540;
  reg  mag_logMagMux_magModule_Queue_1__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_541;
  wire  mag_logMagMux_magModule_Queue_1__T_2; // @[Decoupled.scala 214:41]
  wire  mag_logMagMux_magModule_Queue_1__T_3; // @[Decoupled.scala 215:36]
  wire  mag_logMagMux_magModule_Queue_1__T_4; // @[Decoupled.scala 215:33]
  wire  mag_logMagMux_magModule_Queue_1__T_5; // @[Decoupled.scala 216:32]
  wire  mag_logMagMux_magModule_Queue_1__T_6; // @[Decoupled.scala 40:37]
  wire  mag_logMagMux_magModule_Queue_1__T_8; // @[Decoupled.scala 40:37]
  wire [1:0] mag_logMagMux_magModule_Queue_1__T_12; // @[Counter.scala 39:22]
  wire [1:0] mag_logMagMux_magModule_Queue_1__T_14; // @[Counter.scala 39:22]
  wire  mag_logMagMux_magModule_Queue_1__T_15; // @[Decoupled.scala 227:16]
  wire  mag_logMagMux_magModule__T_2; // @[FixedPointTypeClass.scala 224:24]
  wire [15:0] mag_logMagMux_magModule__T_5; // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] mag_logMagMux_magModule_absInReal; // @[FixedPointTypeClass.scala 247:8]
  wire  mag_logMagMux_magModule__T_6; // @[FixedPointTypeClass.scala 224:24]
  wire [15:0] mag_logMagMux_magModule__T_9; // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] mag_logMagMux_magModule_absInImag; // @[FixedPointTypeClass.scala 247:8]
  wire  mag_logMagMux_magModule__T_10; // @[FixedPointTypeClass.scala 55:59]
  wire [15:0] mag_logMagMux_magModule_u; // @[Order.scala 56:31]
  wire  mag_logMagMux_magModule__T_11; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] mag_logMagMux_magModule_v; // @[Order.scala 55:31]
  wire [12:0] mag_logMagMux_magModule__T_12; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] mag_logMagMux_magModule__GEN_16; // @[FixedPointTypeClass.scala 24:22]
  reg [16:0] mag_logMagMux_magModule__T_14; // @[Reg.scala 15:16]
  reg [31:0] _RAND_542;
  reg [16:0] mag_logMagMux_magModule_jplMagOp1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_543;
  wire [12:0] mag_logMagMux_magModule__T_15; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] mag_logMagMux_magModule__GEN_17; // @[FixedPointTypeClass.scala 33:22]
  reg [16:0] mag_logMagMux_magModule_tmpOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_544;
  reg [14:0] mag_logMagMux_magModule__T_18; // @[Reg.scala 15:16]
  reg [31:0] _RAND_545;
  wire [16:0] mag_logMagMux_magModule__GEN_18; // @[FixedPointTypeClass.scala 24:22]
  reg [17:0] mag_logMagMux_magModule_jplMagOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_546;
  reg [31:0] mag_logMagMux_magModule__T_21; // @[Reg.scala 15:16]
  reg [31:0] _RAND_547;
  wire [17:0] mag_logMagMux_magModule__T_22; // @[FixedPointTypeClass.scala 153:43]
  reg [31:0] mag_logMagMux_magModule__T_24; // @[Reg.scala 15:16]
  reg [31:0] _RAND_548;
  wire [17:0] mag_logMagMux_magModule__T_25; // @[FixedPointTypeClass.scala 153:43]
  reg [18:0] mag_logMagMux_magModule_squared_magnitude; // @[Reg.scala 15:16]
  reg [31:0] _RAND_549;
  wire [17:0] mag_logMagMux_magModule__GEN_19; // @[FixedPointTypeClass.scala 55:59]
  wire  mag_logMagMux_magModule__T_33; // @[FixedPointTypeClass.scala 55:59]
  wire [17:0] mag_logMagMux_magModule_jplMag; // @[Order.scala 56:31]
  reg [1:0] mag_logMagMux_magModule__T_34; // @[Reg.scala 15:16]
  reg [31:0] _RAND_550;
  reg [1:0] mag_logMagMux_magModule__T_35; // @[Reg.scala 15:16]
  reg [31:0] _RAND_551;
  wire  mag_logMagMux_magModule__T_38; // @[Mux.scala 68:19]
  wire [18:0] mag_logMagMux_magModule__T_39; // @[Mux.scala 68:16]
  reg [1:0] mag_logMagMux_magModule_queueCounter; // @[Skid.scala 27:31]
  reg [31:0] _RAND_552;
  wire  mag_logMagMux_magModule__T_48; // @[Skid.scala 35:31]
  wire  mag_logMagMux_magModule__T_49; // @[Skid.scala 35:68]
  wire  mag_logMagMux_magModule__T_50; // @[Skid.scala 35:89]
  wire  mag_logMagMux_magModule_skidInData_ready; // @[Skid.scala 35:51]
  wire  mag_logMagMux_magModule__T_40; // @[Decoupled.scala 40:37]
  wire [1:0] mag_logMagMux_magModule__GEN_20; // @[Skid.scala 28:34]
  wire [2:0] mag_logMagMux_magModule__T_41; // @[Skid.scala 28:34]
  wire  mag_logMagMux_magModule__T_42; // @[Decoupled.scala 40:37]
  wire [2:0] mag_logMagMux_magModule__GEN_21; // @[Skid.scala 28:47]
  wire [3:0] mag_logMagMux_magModule__T_43; // @[Skid.scala 28:47]
  reg  mag_logMagMux_magModule__T_46; // @[Reg.scala 27:20]
  reg [31:0] _RAND_553;
  reg  mag_logMagMux_magModule__T_47; // @[Reg.scala 27:20]
  reg [31:0] _RAND_554;
  wire  mag_logMagMux_magModule__T_54; // @[Decoupled.scala 40:37]
  reg  mag_logMagMux_magModule__T_56; // @[Reg.scala 15:16]
  reg [31:0] _RAND_555;
  reg  mag_logMagMux_magModule__T_57; // @[Reg.scala 15:16]
  reg [31:0] _RAND_556;
  reg [1:0] mag_logMagMux_magModule_queueCounter_1; // @[Skid.scala 27:31]
  reg [31:0] _RAND_557;
  wire  mag_logMagMux_magModule__T_66; // @[Skid.scala 35:31]
  wire  mag_logMagMux_magModule__T_67; // @[Skid.scala 35:68]
  wire  mag_logMagMux_magModule__T_68; // @[Skid.scala 35:89]
  wire  mag_logMagMux_magModule__T_69; // @[Skid.scala 35:51]
  wire  mag_logMagMux_magModule__T_58; // @[Decoupled.scala 40:37]
  wire [1:0] mag_logMagMux_magModule__GEN_22; // @[Skid.scala 28:34]
  wire [2:0] mag_logMagMux_magModule__T_59; // @[Skid.scala 28:34]
  wire  mag_logMagMux_magModule__T_53_valid; // @[LogMagMuxTypes.scala 220:27 Skid.scala 37:15]
  wire  mag_logMagMux_magModule__T_60; // @[Decoupled.scala 40:37]
  wire [2:0] mag_logMagMux_magModule__GEN_23; // @[Skid.scala 28:47]
  wire [3:0] mag_logMagMux_magModule__T_61; // @[Skid.scala 28:47]
  reg  mag_logMagMux_magModule__T_64; // @[Reg.scala 27:20]
  reg [31:0] _RAND_558;
  reg  mag_logMagMux_magModule__T_65; // @[Reg.scala 27:20]
  reg [31:0] _RAND_559;
  wire  mag_Queue_clock;
  wire  mag_Queue_reset;
  wire  mag_Queue_io_enq_ready;
  wire  mag_Queue_io_enq_valid;
  wire  mag_Queue_io_enq_bits_read;
  wire [31:0] mag_Queue_io_enq_bits_data;
  wire  mag_Queue_io_enq_bits_extra;
  wire  mag_Queue_io_deq_ready;
  wire  mag_Queue_io_deq_valid;
  wire  mag_Queue_io_deq_bits_read;
  wire [31:0] mag_Queue_io_deq_bits_data;
  wire  mag_Queue_io_deq_bits_extra;
  reg  mag_Queue__T_read [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_560;
  wire  mag_Queue__T_read__T_18_data; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_read__T_18_addr; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_read__T_10_data; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_read__T_10_addr; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_read__T_10_mask; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_read__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] mag_Queue__T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_561;
  wire [31:0] mag_Queue__T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] mag_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  mag_Queue__T_extra [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_562;
  wire  mag_Queue__T_extra__T_18_data; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_extra__T_18_addr; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_extra__T_10_data; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_extra__T_10_addr; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_extra__T_10_mask; // @[Decoupled.scala 209:24]
  wire  mag_Queue__T_extra__T_10_en; // @[Decoupled.scala 209:24]
  reg  mag_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_563;
  reg  mag_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_564;
  reg  mag_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_565;
  wire  mag_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  mag_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  mag_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  mag_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  mag_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  mag_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  mag_Queue__T_12; // @[Counter.scala 39:22]
  wire  mag_Queue__T_14; // @[Counter.scala 39:22]
  wire  mag_Queue__T_15; // @[Decoupled.scala 227:16]
  reg  mag_selReg; // @[LogMagMuxDspBlock.scala 75:25]
  reg [31:0] _RAND_566;
  wire  mag__T_2; // @[RegisterRouter.scala 40:39]
  wire  mag__T_3; // @[RegisterRouter.scala 40:26]
  wire  mag__T_4; // @[RegisterRouter.scala 42:29]
  wire  mag__T_47_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] mag__T_11; // @[RegisterRouter.scala 48:19]
  wire [27:0] mag__T_45; // @[RegisterRouter.scala 52:27]
  wire [5:0] mag__T_1_bits_index; // @[RegisterRouter.scala 37:18 RegisterRouter.scala 52:19]
  wire  mag__T_53; // @[RegisterRouter.scala 59:16]
  wire  mag__T_5; // @[RegisterRouter.scala 42:26]
  wire  mag__T_13; // @[OneHot.scala 64:49]
  wire [1:0] mag__T_14; // @[OneHot.scala 65:12]
  wire [1:0] mag__T_16; // @[Misc.scala 200:81]
  wire  mag__T_17; // @[Misc.scala 204:21]
  wire  mag__T_18; // @[Misc.scala 207:26]
  wire  mag__T_19; // @[Misc.scala 208:26]
  wire  mag__T_20; // @[Misc.scala 209:20]
  wire  mag__T_22; // @[Misc.scala 213:38]
  wire  mag__T_23; // @[Misc.scala 213:29]
  wire  mag__T_25; // @[Misc.scala 213:38]
  wire  mag__T_26; // @[Misc.scala 213:29]
  wire  mag__T_27; // @[Misc.scala 207:26]
  wire  mag__T_28; // @[Misc.scala 208:26]
  wire  mag__T_29; // @[Misc.scala 209:20]
  wire  mag__T_30; // @[Misc.scala 212:27]
  wire  mag__T_31; // @[Misc.scala 213:38]
  wire  mag__T_32; // @[Misc.scala 213:29]
  wire  mag__T_33; // @[Misc.scala 212:27]
  wire  mag__T_34; // @[Misc.scala 213:38]
  wire  mag__T_35; // @[Misc.scala 213:29]
  wire  mag__T_36; // @[Misc.scala 212:27]
  wire  mag__T_37; // @[Misc.scala 213:38]
  wire  mag__T_38; // @[Misc.scala 213:29]
  wire  mag__T_39; // @[Misc.scala 212:27]
  wire  mag__T_40; // @[Misc.scala 213:38]
  wire  mag__T_41; // @[Misc.scala 213:29]
  wire [3:0] mag__T_44; // @[Cat.scala 29:58]
  wire [3:0] mag__T_46; // @[RegisterRouter.scala 54:25]
  wire  mag__T_58; // @[Bitwise.scala 26:51]
  wire  mag__T_59; // @[Bitwise.scala 26:51]
  wire  mag__T_60; // @[Bitwise.scala 26:51]
  wire  mag__T_61; // @[Bitwise.scala 26:51]
  wire [7:0] mag__T_63; // @[Bitwise.scala 72:12]
  wire [7:0] mag__T_65; // @[Bitwise.scala 72:12]
  wire [7:0] mag__T_67; // @[Bitwise.scala 72:12]
  wire [7:0] mag__T_69; // @[Bitwise.scala 72:12]
  wire [31:0] mag__T_72; // @[Cat.scala 29:58]
  wire  mag__T_88; // @[RegisterRouter.scala 59:16]
  wire  mag__T_117; // @[RegisterRouter.scala 59:16]
  wire  mag__T_129; // @[RegisterRouter.scala 59:16]
  wire  mag__T_132; // @[RegisterRouter.scala 59:16]
  wire  mag__T_98; // @[RegisterRouter.scala 59:16]
  wire  mag__T_100; // @[RegisterRouter.scala 59:16]
  wire  mag__T_171; // @[RegisterRouter.scala 59:16]
  wire  mag__T_172_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  mag__T_172_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  mag__T_175; // @[RegisterRouter.scala 65:29]
  wire  cfar_clock;
  wire  cfar_reset;
  wire  cfar_auto_mem_in_aw_ready;
  wire  cfar_auto_mem_in_aw_valid;
  wire  cfar_auto_mem_in_aw_bits_id;
  wire [29:0] cfar_auto_mem_in_aw_bits_addr;
  wire  cfar_auto_mem_in_w_ready;
  wire  cfar_auto_mem_in_w_valid;
  wire [31:0] cfar_auto_mem_in_w_bits_data;
  wire [3:0] cfar_auto_mem_in_w_bits_strb;
  wire  cfar_auto_mem_in_b_ready;
  wire  cfar_auto_mem_in_b_valid;
  wire  cfar_auto_mem_in_b_bits_id;
  wire  cfar_auto_mem_in_ar_ready;
  wire  cfar_auto_mem_in_ar_valid;
  wire  cfar_auto_mem_in_ar_bits_id;
  wire [29:0] cfar_auto_mem_in_ar_bits_addr;
  wire [2:0] cfar_auto_mem_in_ar_bits_size;
  wire  cfar_auto_mem_in_r_ready;
  wire  cfar_auto_mem_in_r_valid;
  wire  cfar_auto_mem_in_r_bits_id;
  wire [31:0] cfar_auto_mem_in_r_bits_data;
  wire  cfar_auto_master_out_ready;
  wire  cfar_auto_master_out_valid;
  wire [47:0] cfar_auto_master_out_bits_data;
  wire  cfar_auto_master_out_bits_last;
  wire  cfar_auto_slave_in_ready;
  wire  cfar_auto_slave_in_valid;
  wire [15:0] cfar_auto_slave_in_bits_data;
  wire  cfar_auto_slave_in_bits_last;
  wire  cfar_cfar_clock;
  wire  cfar_cfar_reset;
  wire  cfar_cfar_io_in_ready;
  wire  cfar_cfar_io_in_valid;
  wire [15:0] cfar_cfar_io_in_bits;
  wire  cfar_cfar_io_lastIn;
  wire [9:0] cfar_cfar_io_fftWin;
  wire [15:0] cfar_cfar_io_thresholdScaler;
  wire [2:0] cfar_cfar_io_divSum;
  wire  cfar_cfar_io_peakGrouping;
  wire [1:0] cfar_cfar_io_cfarMode;
  wire [6:0] cfar_cfar_io_windowCells;
  wire [3:0] cfar_cfar_io_guardCells;
  wire  cfar_cfar_io_out_ready;
  wire  cfar_cfar_io_out_valid;
  wire  cfar_cfar_io_out_bits_peak;
  wire [15:0] cfar_cfar_io_out_bits_cut;
  wire [15:0] cfar_cfar_io_out_bits_threshold;
  wire  cfar_cfar_io_lastOut;
  wire [8:0] cfar_cfar_io_fftBin;
  wire  cfar_cfar_cfarCore_clock;
  wire  cfar_cfar_cfarCore_reset;
  wire  cfar_cfar_cfarCore_io_in_ready;
  wire  cfar_cfar_cfarCore_io_in_valid;
  wire [15:0] cfar_cfar_cfarCore_io_in_bits;
  wire  cfar_cfar_cfarCore_io_lastIn;
  wire [9:0] cfar_cfar_cfarCore_io_fftWin;
  wire [15:0] cfar_cfar_cfarCore_io_thresholdScaler;
  wire [2:0] cfar_cfar_cfarCore_io_divSum;
  wire  cfar_cfar_cfarCore_io_peakGrouping;
  wire [1:0] cfar_cfar_cfarCore_io_cfarMode;
  wire [6:0] cfar_cfar_cfarCore_io_windowCells;
  wire [3:0] cfar_cfar_cfarCore_io_guardCells;
  wire  cfar_cfar_cfarCore_io_out_ready;
  wire  cfar_cfar_cfarCore_io_out_valid;
  wire  cfar_cfar_cfarCore_io_out_bits_peak;
  wire [15:0] cfar_cfar_cfarCore_io_out_bits_cut;
  wire [15:0] cfar_cfar_cfarCore_io_out_bits_threshold;
  wire  cfar_cfar_cfarCore_io_lastOut;
  wire [8:0] cfar_cfar_cfarCore_io_fftBin;
  wire  cfar_cfar_cfarCore_laggWindow_clock;
  wire  cfar_cfar_cfarCore_laggWindow_reset;
  wire [6:0] cfar_cfar_cfarCore_laggWindow_io_depth;
  wire  cfar_cfar_cfarCore_laggWindow_io_in_ready;
  wire  cfar_cfar_cfarCore_laggWindow_io_in_valid;
  wire [15:0] cfar_cfar_cfarCore_laggWindow_io_in_bits;
  wire  cfar_cfar_cfarCore_laggWindow_io_lastIn;
  wire  cfar_cfar_cfarCore_laggWindow_io_out_ready;
  wire  cfar_cfar_cfarCore_laggWindow_io_out_valid;
  wire [15:0] cfar_cfar_cfarCore_laggWindow_io_out_bits;
  wire  cfar_cfar_cfarCore_laggWindow_io_lastOut;
  wire  cfar_cfar_cfarCore_laggWindow_io_memFull;
  reg [15:0] cfar_cfar_cfarCore_laggWindow_mem [0:63]; // @[CFARUtils.scala 505:26]
  reg [31:0] _RAND_567;
  wire [15:0] cfar_cfar_cfarCore_laggWindow_mem__T_423_data; // @[CFARUtils.scala 505:26]
  wire [5:0] cfar_cfar_cfarCore_laggWindow_mem__T_423_addr; // @[CFARUtils.scala 505:26]
  wire [15:0] cfar_cfar_cfarCore_laggWindow_mem__T_418_data; // @[CFARUtils.scala 505:26]
  wire [5:0] cfar_cfar_cfarCore_laggWindow_mem__T_418_addr; // @[CFARUtils.scala 505:26]
  wire  cfar_cfar_cfarCore_laggWindow_mem__T_418_mask; // @[CFARUtils.scala 505:26]
  wire  cfar_cfar_cfarCore_laggWindow_mem__T_418_en; // @[CFARUtils.scala 505:26]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue_clock;
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue_reset;
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_ready;
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_valid;
  wire [15:0] cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_bits;
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_ready;
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_valid;
  wire [15:0] cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_bits;
  reg [15:0] cfar_cfar_cfarCore_laggWindow_outputQueue__T [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_568;
  wire [15:0] cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_14_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_14_addr; // @[Decoupled.scala 209:24]
  wire [15:0] cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_en; // @[Decoupled.scala 209:24]
  reg  cfar_cfar_cfarCore_laggWindow_outputQueue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_569;
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T_3; // @[Decoupled.scala 215:36]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T_6; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T_8; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_7; // @[Decoupled.scala 240:27]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_10; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_9; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T_11; // @[Decoupled.scala 227:16]
  wire  cfar_cfar_cfarCore_laggWindow_outputQueue__T_12; // @[Decoupled.scala 231:19]
  reg [5:0] cfar_cfar_cfarCore_laggWindow_writeIdxReg; // @[CFARUtils.scala 508:30]
  reg [31:0] _RAND_570;
  reg  cfar_cfar_cfarCore_laggWindow_last; // @[CFARUtils.scala 509:30]
  reg [31:0] _RAND_571;
  reg  cfar_cfar_cfarCore_laggWindow_initialInDone; // @[CFARUtils.scala 510:30]
  reg [31:0] _RAND_572;
  wire  cfar_cfar_cfarCore_laggWindow__T; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_1; // @[CFARUtils.scala 511:45]
  wire  cfar_cfar_cfarCore_laggWindow_en; // @[CFARUtils.scala 511:36]
  reg  cfar_cfar_cfarCore_laggWindow_validPrev; // @[CFARUtils.scala 514:26]
  reg [31:0] _RAND_573;
  wire [5:0] cfar_cfar_cfarCore_laggWindow__T_3; // @[CFARUtils.scala 515:21]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__GEN_140; // @[CFARUtils.scala 515:27]
  wire  cfar_cfar_cfarCore_laggWindow__T_4; // @[CFARUtils.scala 515:27]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__GEN_141; // @[CFARUtils.scala 516:28]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__T_6; // @[CFARUtils.scala 516:28]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__T_8; // @[CFARUtils.scala 516:39]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__T_10; // @[CFARUtils.scala 518:27]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__T_12; // @[CFARUtils.scala 518:41]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__T_14; // @[CFARUtils.scala 518:47]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__GEN_0; // @[CFARUtils.scala 515:40]
  wire [6:0] cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 528:34]
  wire  cfar_cfar_cfarCore_laggWindow__T_17; // @[CFARUtils.scala 528:21]
  wire  cfar_cfar_cfarCore_laggWindow__T_19; // @[CFARUtils.scala 528:40]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_1; // @[CFARUtils.scala 528:57]
  wire  cfar_cfar_cfarCore_laggWindow_fireLastIn; // @[CFARUtils.scala 531:30]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_2; // @[CFARUtils.scala 533:21]
  wire  cfar_cfar_cfarCore_laggWindow__T_21; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_22; // @[CFARUtils.scala 330:18]
  wire  cfar_cfar_cfarCore_laggWindow__T_24; // @[CFARUtils.scala 330:11]
  wire  cfar_cfar_cfarCore_laggWindow__T_25; // @[CFARUtils.scala 330:11]
  wire  cfar_cfar_cfarCore_laggWindow__T_33; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_37; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_41; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_45; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_49; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_53; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_57; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_61; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_65; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_69; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_73; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_77; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_81; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_85; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_89; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_93; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_97; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_101; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_105; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_109; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_113; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_117; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_121; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_125; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_129; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_133; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_137; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_141; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_145; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_149; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_153; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_157; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_161; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_165; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_169; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_173; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_177; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_181; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_185; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_189; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_193; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_197; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_201; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_205; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_209; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_213; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_217; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_221; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_225; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_229; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_233; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_237; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_241; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_245; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_249; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_253; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_257; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_261; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_265; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_269; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_273; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_277; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_281; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_laggWindow__T_284; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_285; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_286; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_287; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_288; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_289; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_290; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_291; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_292; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_293; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_294; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_295; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_296; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_297; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_298; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_299; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_300; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_301; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_302; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_303; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_304; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_305; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_306; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_307; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_308; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_309; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_310; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_311; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_312; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_313; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_314; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_315; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_316; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_317; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_318; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_319; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_320; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_321; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_322; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_323; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_324; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_325; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_326; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_327; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_328; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_329; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_330; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_331; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_332; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_333; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_334; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_335; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_336; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_337; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_338; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_339; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_340; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_341; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_342; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_343; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_344; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_345; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggWindow__T_346; // @[CFARUtils.scala 319:37]
  reg  cfar_cfar_cfarCore_laggWindow__T_348; // @[Reg.scala 27:20]
  reg [31:0] _RAND_574;
  reg  cfar_cfar_cfarCore_laggWindow__T_349; // @[Reg.scala 27:20]
  reg [31:0] _RAND_575;
  reg  cfar_cfar_cfarCore_laggWindow__T_350; // @[Reg.scala 27:20]
  reg [31:0] _RAND_576;
  reg  cfar_cfar_cfarCore_laggWindow__T_351; // @[Reg.scala 27:20]
  reg [31:0] _RAND_577;
  reg  cfar_cfar_cfarCore_laggWindow__T_352; // @[Reg.scala 27:20]
  reg [31:0] _RAND_578;
  reg  cfar_cfar_cfarCore_laggWindow__T_353; // @[Reg.scala 27:20]
  reg [31:0] _RAND_579;
  reg  cfar_cfar_cfarCore_laggWindow__T_354; // @[Reg.scala 27:20]
  reg [31:0] _RAND_580;
  reg  cfar_cfar_cfarCore_laggWindow__T_355; // @[Reg.scala 27:20]
  reg [31:0] _RAND_581;
  reg  cfar_cfar_cfarCore_laggWindow__T_356; // @[Reg.scala 27:20]
  reg [31:0] _RAND_582;
  reg  cfar_cfar_cfarCore_laggWindow__T_357; // @[Reg.scala 27:20]
  reg [31:0] _RAND_583;
  reg  cfar_cfar_cfarCore_laggWindow__T_358; // @[Reg.scala 27:20]
  reg [31:0] _RAND_584;
  reg  cfar_cfar_cfarCore_laggWindow__T_359; // @[Reg.scala 27:20]
  reg [31:0] _RAND_585;
  reg  cfar_cfar_cfarCore_laggWindow__T_360; // @[Reg.scala 27:20]
  reg [31:0] _RAND_586;
  reg  cfar_cfar_cfarCore_laggWindow__T_361; // @[Reg.scala 27:20]
  reg [31:0] _RAND_587;
  reg  cfar_cfar_cfarCore_laggWindow__T_362; // @[Reg.scala 27:20]
  reg [31:0] _RAND_588;
  reg  cfar_cfar_cfarCore_laggWindow__T_363; // @[Reg.scala 27:20]
  reg [31:0] _RAND_589;
  reg  cfar_cfar_cfarCore_laggWindow__T_364; // @[Reg.scala 27:20]
  reg [31:0] _RAND_590;
  reg  cfar_cfar_cfarCore_laggWindow__T_365; // @[Reg.scala 27:20]
  reg [31:0] _RAND_591;
  reg  cfar_cfar_cfarCore_laggWindow__T_366; // @[Reg.scala 27:20]
  reg [31:0] _RAND_592;
  reg  cfar_cfar_cfarCore_laggWindow__T_367; // @[Reg.scala 27:20]
  reg [31:0] _RAND_593;
  reg  cfar_cfar_cfarCore_laggWindow__T_368; // @[Reg.scala 27:20]
  reg [31:0] _RAND_594;
  reg  cfar_cfar_cfarCore_laggWindow__T_369; // @[Reg.scala 27:20]
  reg [31:0] _RAND_595;
  reg  cfar_cfar_cfarCore_laggWindow__T_370; // @[Reg.scala 27:20]
  reg [31:0] _RAND_596;
  reg  cfar_cfar_cfarCore_laggWindow__T_371; // @[Reg.scala 27:20]
  reg [31:0] _RAND_597;
  reg  cfar_cfar_cfarCore_laggWindow__T_372; // @[Reg.scala 27:20]
  reg [31:0] _RAND_598;
  reg  cfar_cfar_cfarCore_laggWindow__T_373; // @[Reg.scala 27:20]
  reg [31:0] _RAND_599;
  reg  cfar_cfar_cfarCore_laggWindow__T_374; // @[Reg.scala 27:20]
  reg [31:0] _RAND_600;
  reg  cfar_cfar_cfarCore_laggWindow__T_375; // @[Reg.scala 27:20]
  reg [31:0] _RAND_601;
  reg  cfar_cfar_cfarCore_laggWindow__T_376; // @[Reg.scala 27:20]
  reg [31:0] _RAND_602;
  reg  cfar_cfar_cfarCore_laggWindow__T_377; // @[Reg.scala 27:20]
  reg [31:0] _RAND_603;
  reg  cfar_cfar_cfarCore_laggWindow__T_378; // @[Reg.scala 27:20]
  reg [31:0] _RAND_604;
  reg  cfar_cfar_cfarCore_laggWindow__T_379; // @[Reg.scala 27:20]
  reg [31:0] _RAND_605;
  reg  cfar_cfar_cfarCore_laggWindow__T_380; // @[Reg.scala 27:20]
  reg [31:0] _RAND_606;
  reg  cfar_cfar_cfarCore_laggWindow__T_381; // @[Reg.scala 27:20]
  reg [31:0] _RAND_607;
  reg  cfar_cfar_cfarCore_laggWindow__T_382; // @[Reg.scala 27:20]
  reg [31:0] _RAND_608;
  reg  cfar_cfar_cfarCore_laggWindow__T_383; // @[Reg.scala 27:20]
  reg [31:0] _RAND_609;
  reg  cfar_cfar_cfarCore_laggWindow__T_384; // @[Reg.scala 27:20]
  reg [31:0] _RAND_610;
  reg  cfar_cfar_cfarCore_laggWindow__T_385; // @[Reg.scala 27:20]
  reg [31:0] _RAND_611;
  reg  cfar_cfar_cfarCore_laggWindow__T_386; // @[Reg.scala 27:20]
  reg [31:0] _RAND_612;
  reg  cfar_cfar_cfarCore_laggWindow__T_387; // @[Reg.scala 27:20]
  reg [31:0] _RAND_613;
  reg  cfar_cfar_cfarCore_laggWindow__T_388; // @[Reg.scala 27:20]
  reg [31:0] _RAND_614;
  reg  cfar_cfar_cfarCore_laggWindow__T_389; // @[Reg.scala 27:20]
  reg [31:0] _RAND_615;
  reg  cfar_cfar_cfarCore_laggWindow__T_390; // @[Reg.scala 27:20]
  reg [31:0] _RAND_616;
  reg  cfar_cfar_cfarCore_laggWindow__T_391; // @[Reg.scala 27:20]
  reg [31:0] _RAND_617;
  reg  cfar_cfar_cfarCore_laggWindow__T_392; // @[Reg.scala 27:20]
  reg [31:0] _RAND_618;
  reg  cfar_cfar_cfarCore_laggWindow__T_393; // @[Reg.scala 27:20]
  reg [31:0] _RAND_619;
  reg  cfar_cfar_cfarCore_laggWindow__T_394; // @[Reg.scala 27:20]
  reg [31:0] _RAND_620;
  reg  cfar_cfar_cfarCore_laggWindow__T_395; // @[Reg.scala 27:20]
  reg [31:0] _RAND_621;
  reg  cfar_cfar_cfarCore_laggWindow__T_396; // @[Reg.scala 27:20]
  reg [31:0] _RAND_622;
  reg  cfar_cfar_cfarCore_laggWindow__T_397; // @[Reg.scala 27:20]
  reg [31:0] _RAND_623;
  reg  cfar_cfar_cfarCore_laggWindow__T_398; // @[Reg.scala 27:20]
  reg [31:0] _RAND_624;
  reg  cfar_cfar_cfarCore_laggWindow__T_399; // @[Reg.scala 27:20]
  reg [31:0] _RAND_625;
  reg  cfar_cfar_cfarCore_laggWindow__T_400; // @[Reg.scala 27:20]
  reg [31:0] _RAND_626;
  reg  cfar_cfar_cfarCore_laggWindow__T_401; // @[Reg.scala 27:20]
  reg [31:0] _RAND_627;
  reg  cfar_cfar_cfarCore_laggWindow__T_402; // @[Reg.scala 27:20]
  reg [31:0] _RAND_628;
  reg  cfar_cfar_cfarCore_laggWindow__T_403; // @[Reg.scala 27:20]
  reg [31:0] _RAND_629;
  reg  cfar_cfar_cfarCore_laggWindow__T_404; // @[Reg.scala 27:20]
  reg [31:0] _RAND_630;
  reg  cfar_cfar_cfarCore_laggWindow__T_405; // @[Reg.scala 27:20]
  reg [31:0] _RAND_631;
  reg  cfar_cfar_cfarCore_laggWindow__T_406; // @[Reg.scala 27:20]
  reg [31:0] _RAND_632;
  reg  cfar_cfar_cfarCore_laggWindow__T_407; // @[Reg.scala 27:20]
  reg [31:0] _RAND_633;
  reg  cfar_cfar_cfarCore_laggWindow__T_408; // @[Reg.scala 27:20]
  reg [31:0] _RAND_634;
  reg  cfar_cfar_cfarCore_laggWindow__T_409; // @[Reg.scala 27:20]
  reg [31:0] _RAND_635;
  reg  cfar_cfar_cfarCore_laggWindow__T_410; // @[Reg.scala 27:20]
  reg [31:0] _RAND_636;
  reg  cfar_cfar_cfarCore_laggWindow__T_411; // @[Reg.scala 27:20]
  reg [31:0] _RAND_637;
  wire [5:0] cfar_cfar_cfarCore_laggWindow__T_414;
  wire  cfar_cfar_cfarCore_laggWindow__GEN_68; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_69; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_70; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_71; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_72; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_73; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_74; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_75; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_76; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_77; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_78; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_79; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_80; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_81; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_82; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_83; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_84; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_85; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_86; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_87; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_88; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_89; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_90; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_91; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_92; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_93; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_94; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_95; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_96; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_97; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_98; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_99; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_100; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_101; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_102; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_103; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_104; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_105; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_106; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_107; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_108; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_109; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_110; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_111; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_112; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_113; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_114; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_115; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_116; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_117; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_118; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_119; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_120; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_121; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_122; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_123; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_124; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_125; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_126; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_127; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_128; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_129; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__GEN_130; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow_resetAll; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_laggWindow__T_416; // @[CFARUtils.scala 544:15]
  wire  cfar_cfar_cfarCore_laggWindow__T_417; // @[CFARUtils.scala 544:12]
  wire  cfar_cfar_cfarCore_laggWindow__T_419; // @[CFARUtils.scala 546:36]
  reg [15:0] cfar_cfar_cfarCore_laggWindow__T_426; // @[CFARUtils.scala 551:37]
  reg [31:0] _RAND_638;
  wire  cfar_cfar_cfarCore_laggWindow__T_431; // @[CFARUtils.scala 554:42]
  wire  cfar_cfar_cfarCore_laggWindow__T_433; // @[CFARUtils.scala 555:36]
  wire  cfar_cfar_cfarCore_laggWindow__T_437; // @[CFARUtils.scala 559:52]
  wire  cfar_cfar_cfarCore_laggWindow__T_439; // @[CFARUtils.scala 568:33]
  wire  cfar_cfar_cfarCore_laggWindow__T_440; // @[CFARUtils.scala 568:57]
  wire [5:0] cfar_cfar_cfarCore_laggWindow_readIdx; // @[CFARUtils.scala 506:27 CFARUtils.scala 516:13 CFARUtils.scala 518:13]
  wire  cfar_cfar_cfarCore_laggGuard_clock;
  wire  cfar_cfar_cfarCore_laggGuard_reset;
  wire [3:0] cfar_cfar_cfarCore_laggGuard_io_depth;
  wire  cfar_cfar_cfarCore_laggGuard_io_in_ready;
  wire  cfar_cfar_cfarCore_laggGuard_io_in_valid;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_in_bits;
  wire  cfar_cfar_cfarCore_laggGuard_io_lastIn;
  wire  cfar_cfar_cfarCore_laggGuard_io_out_ready;
  wire  cfar_cfar_cfarCore_laggGuard_io_out_valid;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_out_bits;
  wire  cfar_cfar_cfarCore_laggGuard_io_lastOut;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_0;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_1;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_2;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_3;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_4;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_5;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_6;
  wire [15:0] cfar_cfar_cfarCore_laggGuard_io_parallelOut_7;
  reg  cfar_cfar_cfarCore_laggGuard_InitialInDone; // @[CFARUtils.scala 379:30]
  reg [31:0] _RAND_639;
  reg  cfar_cfar_cfarCore_laggGuard_last; // @[CFARUtils.scala 380:21]
  reg [31:0] _RAND_640;
  wire  cfar_cfar_cfarCore_laggGuard__T_1; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_2; // @[CFARUtils.scala 385:34]
  wire  cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 385:25]
  wire  cfar_cfar_cfarCore_laggGuard__T_3; // @[CFARUtils.scala 345:18]
  wire  cfar_cfar_cfarCore_laggGuard__T_5; // @[CFARUtils.scala 345:11]
  wire  cfar_cfar_cfarCore_laggGuard__T_6; // @[CFARUtils.scala 345:11]
  wire [3:0] cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:87]
  wire  cfar_cfar_cfarCore_laggGuard__T_9; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_13; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_14; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_17; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_18; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_21; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_22; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_25; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_26; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_29; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_30; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_33; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_34; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_37; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_laggGuard__T_38; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_39; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_40; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_41; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_42; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_43; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_44; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_45; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_46; // @[CFARUtils.scala 319:37]
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_641;
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_1; // @[Reg.scala 27:20]
  reg [31:0] _RAND_642;
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_2; // @[Reg.scala 27:20]
  reg [31:0] _RAND_643;
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_3; // @[Reg.scala 27:20]
  reg [31:0] _RAND_644;
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_4; // @[Reg.scala 27:20]
  reg [31:0] _RAND_645;
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_5; // @[Reg.scala 27:20]
  reg [31:0] _RAND_646;
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_6; // @[Reg.scala 27:20]
  reg [31:0] _RAND_647;
  reg [15:0] cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_7; // @[Reg.scala 27:20]
  reg [31:0] _RAND_648;
  wire [2:0] cfar_cfar_cfarCore_laggGuard__T_57;
  reg [3:0] cfar_cfar_cfarCore_laggGuard_cntIn; // @[CFARUtils.scala 390:23]
  reg [31:0] _RAND_649;
  wire  cfar_cfar_cfarCore_laggGuard__T_59; // @[CFARUtils.scala 392:19]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_8; // @[CFARUtils.scala 392:36]
  wire [3:0] cfar_cfar_cfarCore_laggGuard__T_62; // @[CFARUtils.scala 397:20]
  wire  cfar_cfar_cfarCore_laggGuard__T_63; // @[CFARUtils.scala 400:18]
  wire  cfar_cfar_cfarCore_laggGuard__T_66; // @[CFARUtils.scala 401:17]
  wire  cfar_cfar_cfarCore_laggGuard__T_68; // @[CFARUtils.scala 401:36]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_10; // @[CFARUtils.scala 401:53]
  wire  cfar_cfar_cfarCore_laggGuard__T_70; // @[CFARUtils.scala 406:36]
  wire  cfar_cfar_cfarCore_laggGuard__T_71; // @[CFARUtils.scala 406:24]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_11; // @[CFARUtils.scala 406:45]
  wire  cfar_cfar_cfarCore_laggGuard__T_73; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_112; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_113; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_114; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_115; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_116; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_117; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_118; // @[CFARUtils.scala 319:37]
  reg  cfar_cfar_cfarCore_laggGuard__T_120; // @[Reg.scala 27:20]
  reg [31:0] _RAND_650;
  reg  cfar_cfar_cfarCore_laggGuard__T_121; // @[Reg.scala 27:20]
  reg [31:0] _RAND_651;
  reg  cfar_cfar_cfarCore_laggGuard__T_122; // @[Reg.scala 27:20]
  reg [31:0] _RAND_652;
  reg  cfar_cfar_cfarCore_laggGuard__T_123; // @[Reg.scala 27:20]
  reg [31:0] _RAND_653;
  reg  cfar_cfar_cfarCore_laggGuard__T_124; // @[Reg.scala 27:20]
  reg [31:0] _RAND_654;
  reg  cfar_cfar_cfarCore_laggGuard__T_125; // @[Reg.scala 27:20]
  reg [31:0] _RAND_655;
  reg  cfar_cfar_cfarCore_laggGuard__T_126; // @[Reg.scala 27:20]
  reg [31:0] _RAND_656;
  reg  cfar_cfar_cfarCore_laggGuard__T_127; // @[Reg.scala 27:20]
  reg [31:0] _RAND_657;
  wire  cfar_cfar_cfarCore_laggGuard__GEN_22; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_23; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_24; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_25; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_26; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_27; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__GEN_28; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__T_132; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_laggGuard__T_134; // @[CFARUtils.scala 420:36]
  wire  cfar_cfar_cfarCore_laggGuard__T_136; // @[CFARUtils.scala 421:36]
  wire  cfar_cfar_cfarCore_laggGuard__T_138; // @[CFARUtils.scala 426:37]
  wire  cfar_cfar_cfarCore_laggGuard__T_141; // @[CFARUtils.scala 426:91]
  wire  cfar_cfar_cfarCore_laggGuard__T_142; // @[CFARUtils.scala 426:75]
  wire [15:0] cfar_cfar_cfarCore_laggGuard__GEN_33; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_laggGuard__GEN_34; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_laggGuard__GEN_35; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_laggGuard__GEN_36; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_laggGuard__GEN_37; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_laggGuard__GEN_38; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_laggGuard__GEN_39; // @[CFARUtils.scala 433:24]
  wire  cfar_cfar_cfarCore_laggGuard__T_151; // @[CFARUtils.scala 436:70]
  wire  cfar_cfar_cfarCore_laggGuard__T_152; // @[CFARUtils.scala 436:94]
  wire  cfar_cfar_cfarCore_laggGuard__T_153; // @[CFARUtils.scala 436:85]
  wire  cfar_cfar_cfarCore_cellUnderTest_clock;
  wire  cfar_cfar_cfarCore_cellUnderTest_reset;
  wire  cfar_cfar_cfarCore_cellUnderTest_io_in_ready;
  wire  cfar_cfar_cfarCore_cellUnderTest_io_in_valid;
  wire [15:0] cfar_cfar_cfarCore_cellUnderTest_io_in_bits;
  wire  cfar_cfar_cfarCore_cellUnderTest_io_lastIn;
  wire  cfar_cfar_cfarCore_cellUnderTest_io_out_ready;
  wire  cfar_cfar_cfarCore_cellUnderTest_io_out_valid;
  wire [15:0] cfar_cfar_cfarCore_cellUnderTest_io_out_bits;
  wire  cfar_cfar_cfarCore_cellUnderTest_io_lastOut;
  reg  cfar_cfar_cfarCore_cellUnderTest_initialInDone; // @[CFARUtils.scala 453:30]
  reg [31:0] _RAND_658;
  reg  cfar_cfar_cfarCore_cellUnderTest_last; // @[CFARUtils.scala 455:21]
  reg [31:0] _RAND_659;
  wire  cfar_cfar_cfarCore_cellUnderTest__T_1; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_cellUnderTest__T_2; // @[CFARUtils.scala 457:25]
  wire  cfar_cfar_cfarCore_cellUnderTest__T_3; // @[CFARUtils.scala 457:22]
  wire  cfar_cfar_cfarCore_cellUnderTest__GEN_0; // @[CFARUtils.scala 457:41]
  wire  cfar_cfar_cfarCore_cellUnderTest__T_5; // @[CFARUtils.scala 461:34]
  wire  cfar_cfar_cfarCore_cellUnderTest_en; // @[CFARUtils.scala 461:25]
  reg [15:0] cfar_cfar_cfarCore_cellUnderTest_cut; // @[Reg.scala 27:20]
  reg [31:0] _RAND_660;
  wire  cfar_cfar_cfarCore_cellUnderTest__T_7; // @[CFARUtils.scala 468:19]
  wire  cfar_cfar_cfarCore_cellUnderTest__GEN_2; // @[CFARUtils.scala 468:36]
  reg  cfar_cfar_cfarCore_cellUnderTest_lastOut; // @[Reg.scala 27:20]
  reg [31:0] _RAND_661;
  wire  cfar_cfar_cfarCore_cellUnderTest__T_9; // @[CFARUtils.scala 475:17]
  wire  cfar_cfar_cfarCore_cellUnderTest__T_11; // @[CFARUtils.scala 480:55]
  wire  cfar_cfar_cfarCore_cellUnderTest__T_12; // @[CFARUtils.scala 480:52]
  wire  cfar_cfar_cfarCore_cellUnderTest__T_14; // @[CFARUtils.scala 483:35]
  wire  cfar_cfar_cfarCore_cellUnderTest__T_15; // @[CFARUtils.scala 483:59]
  wire  cfar_cfar_cfarCore_leadGuard_clock;
  wire  cfar_cfar_cfarCore_leadGuard_reset;
  wire [3:0] cfar_cfar_cfarCore_leadGuard_io_depth;
  wire  cfar_cfar_cfarCore_leadGuard_io_in_ready;
  wire  cfar_cfar_cfarCore_leadGuard_io_in_valid;
  wire [15:0] cfar_cfar_cfarCore_leadGuard_io_in_bits;
  wire  cfar_cfar_cfarCore_leadGuard_io_lastIn;
  wire  cfar_cfar_cfarCore_leadGuard_io_out_ready;
  wire  cfar_cfar_cfarCore_leadGuard_io_out_valid;
  wire [15:0] cfar_cfar_cfarCore_leadGuard_io_out_bits;
  wire  cfar_cfar_cfarCore_leadGuard_io_lastOut;
  reg  cfar_cfar_cfarCore_leadGuard_InitialInDone; // @[CFARUtils.scala 379:30]
  reg [31:0] _RAND_662;
  reg  cfar_cfar_cfarCore_leadGuard_last; // @[CFARUtils.scala 380:21]
  reg [31:0] _RAND_663;
  wire  cfar_cfar_cfarCore_leadGuard__T_1; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_2; // @[CFARUtils.scala 385:34]
  wire  cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 385:25]
  wire  cfar_cfar_cfarCore_leadGuard__T_3; // @[CFARUtils.scala 345:18]
  wire  cfar_cfar_cfarCore_leadGuard__T_5; // @[CFARUtils.scala 345:11]
  wire  cfar_cfar_cfarCore_leadGuard__T_6; // @[CFARUtils.scala 345:11]
  wire [3:0] cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:87]
  wire  cfar_cfar_cfarCore_leadGuard__T_9; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_13; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_14; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_17; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_18; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_21; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_22; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_25; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_26; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_29; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_30; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_33; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_34; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_37; // @[CFARUtils.scala 350:78]
  wire  cfar_cfar_cfarCore_leadGuard__T_38; // @[CFARUtils.scala 350:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_39; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_40; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_41; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_42; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_43; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_44; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_45; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_46; // @[CFARUtils.scala 319:37]
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_664;
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_1; // @[Reg.scala 27:20]
  reg [31:0] _RAND_665;
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_2; // @[Reg.scala 27:20]
  reg [31:0] _RAND_666;
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_3; // @[Reg.scala 27:20]
  reg [31:0] _RAND_667;
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_4; // @[Reg.scala 27:20]
  reg [31:0] _RAND_668;
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_5; // @[Reg.scala 27:20]
  reg [31:0] _RAND_669;
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_6; // @[Reg.scala 27:20]
  reg [31:0] _RAND_670;
  reg [15:0] cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_7; // @[Reg.scala 27:20]
  reg [31:0] _RAND_671;
  wire [2:0] cfar_cfar_cfarCore_leadGuard__T_57;
  reg [3:0] cfar_cfar_cfarCore_leadGuard_cntIn; // @[CFARUtils.scala 390:23]
  reg [31:0] _RAND_672;
  wire  cfar_cfar_cfarCore_leadGuard__T_59; // @[CFARUtils.scala 392:19]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_8; // @[CFARUtils.scala 392:36]
  wire [3:0] cfar_cfar_cfarCore_leadGuard__T_62; // @[CFARUtils.scala 397:20]
  wire  cfar_cfar_cfarCore_leadGuard__T_63; // @[CFARUtils.scala 400:18]
  wire  cfar_cfar_cfarCore_leadGuard__T_66; // @[CFARUtils.scala 401:17]
  wire  cfar_cfar_cfarCore_leadGuard__T_68; // @[CFARUtils.scala 401:36]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_10; // @[CFARUtils.scala 401:53]
  wire  cfar_cfar_cfarCore_leadGuard__T_70; // @[CFARUtils.scala 406:36]
  wire  cfar_cfar_cfarCore_leadGuard__T_71; // @[CFARUtils.scala 406:24]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_11; // @[CFARUtils.scala 406:45]
  wire  cfar_cfar_cfarCore_leadGuard__T_73; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_112; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_113; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_114; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_115; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_116; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_117; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_118; // @[CFARUtils.scala 319:37]
  reg  cfar_cfar_cfarCore_leadGuard__T_120; // @[Reg.scala 27:20]
  reg [31:0] _RAND_673;
  reg  cfar_cfar_cfarCore_leadGuard__T_121; // @[Reg.scala 27:20]
  reg [31:0] _RAND_674;
  reg  cfar_cfar_cfarCore_leadGuard__T_122; // @[Reg.scala 27:20]
  reg [31:0] _RAND_675;
  reg  cfar_cfar_cfarCore_leadGuard__T_123; // @[Reg.scala 27:20]
  reg [31:0] _RAND_676;
  reg  cfar_cfar_cfarCore_leadGuard__T_124; // @[Reg.scala 27:20]
  reg [31:0] _RAND_677;
  reg  cfar_cfar_cfarCore_leadGuard__T_125; // @[Reg.scala 27:20]
  reg [31:0] _RAND_678;
  reg  cfar_cfar_cfarCore_leadGuard__T_126; // @[Reg.scala 27:20]
  reg [31:0] _RAND_679;
  reg  cfar_cfar_cfarCore_leadGuard__T_127; // @[Reg.scala 27:20]
  reg [31:0] _RAND_680;
  wire  cfar_cfar_cfarCore_leadGuard__GEN_22; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_23; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_24; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_25; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_26; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_27; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__GEN_28; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__T_132; // @[CFARUtils.scala 414:17]
  wire  cfar_cfar_cfarCore_leadGuard__T_134; // @[CFARUtils.scala 420:36]
  wire  cfar_cfar_cfarCore_leadGuard__T_136; // @[CFARUtils.scala 421:36]
  wire  cfar_cfar_cfarCore_leadGuard__T_138; // @[CFARUtils.scala 426:37]
  wire  cfar_cfar_cfarCore_leadGuard__T_141; // @[CFARUtils.scala 426:91]
  wire  cfar_cfar_cfarCore_leadGuard__T_142; // @[CFARUtils.scala 426:75]
  wire [15:0] cfar_cfar_cfarCore_leadGuard__GEN_33; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_leadGuard__GEN_34; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_leadGuard__GEN_35; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_leadGuard__GEN_36; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_leadGuard__GEN_37; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_leadGuard__GEN_38; // @[CFARUtils.scala 433:24]
  wire [15:0] cfar_cfar_cfarCore_leadGuard__GEN_39; // @[CFARUtils.scala 433:24]
  wire  cfar_cfar_cfarCore_leadGuard__T_151; // @[CFARUtils.scala 436:70]
  wire  cfar_cfar_cfarCore_leadGuard__T_152; // @[CFARUtils.scala 436:94]
  wire  cfar_cfar_cfarCore_leadGuard__T_153; // @[CFARUtils.scala 436:85]
  wire  cfar_cfar_cfarCore_leadWindow_clock;
  wire  cfar_cfar_cfarCore_leadWindow_reset;
  wire [6:0] cfar_cfar_cfarCore_leadWindow_io_depth;
  wire  cfar_cfar_cfarCore_leadWindow_io_in_ready;
  wire  cfar_cfar_cfarCore_leadWindow_io_in_valid;
  wire [15:0] cfar_cfar_cfarCore_leadWindow_io_in_bits;
  wire  cfar_cfar_cfarCore_leadWindow_io_lastIn;
  wire  cfar_cfar_cfarCore_leadWindow_io_out_ready;
  wire  cfar_cfar_cfarCore_leadWindow_io_out_valid;
  wire [15:0] cfar_cfar_cfarCore_leadWindow_io_out_bits;
  wire  cfar_cfar_cfarCore_leadWindow_io_memFull;
  wire  cfar_cfar_cfarCore_leadWindow_io_memEmpty;
  reg [15:0] cfar_cfar_cfarCore_leadWindow_mem [0:63]; // @[CFARUtils.scala 505:26]
  reg [31:0] _RAND_681;
  wire [15:0] cfar_cfar_cfarCore_leadWindow_mem__T_423_data; // @[CFARUtils.scala 505:26]
  wire [5:0] cfar_cfar_cfarCore_leadWindow_mem__T_423_addr; // @[CFARUtils.scala 505:26]
  wire [15:0] cfar_cfar_cfarCore_leadWindow_mem__T_418_data; // @[CFARUtils.scala 505:26]
  wire [5:0] cfar_cfar_cfarCore_leadWindow_mem__T_418_addr; // @[CFARUtils.scala 505:26]
  wire  cfar_cfar_cfarCore_leadWindow_mem__T_418_mask; // @[CFARUtils.scala 505:26]
  wire  cfar_cfar_cfarCore_leadWindow_mem__T_418_en; // @[CFARUtils.scala 505:26]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue_clock;
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue_reset;
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_ready;
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_valid;
  wire [15:0] cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_bits;
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_ready;
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_valid;
  wire [15:0] cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_bits;
  reg [15:0] cfar_cfar_cfarCore_leadWindow_outputQueue__T [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_682;
  wire [15:0] cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_14_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_14_addr; // @[Decoupled.scala 209:24]
  wire [15:0] cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_en; // @[Decoupled.scala 209:24]
  reg  cfar_cfar_cfarCore_leadWindow_outputQueue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_683;
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T_3; // @[Decoupled.scala 215:36]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T_6; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T_8; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_7; // @[Decoupled.scala 240:27]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_10; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_9; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T_11; // @[Decoupled.scala 227:16]
  wire  cfar_cfar_cfarCore_leadWindow_outputQueue__T_12; // @[Decoupled.scala 231:19]
  reg [5:0] cfar_cfar_cfarCore_leadWindow_writeIdxReg; // @[CFARUtils.scala 508:30]
  reg [31:0] _RAND_684;
  reg  cfar_cfar_cfarCore_leadWindow_last; // @[CFARUtils.scala 509:30]
  reg [31:0] _RAND_685;
  reg  cfar_cfar_cfarCore_leadWindow_initialInDone; // @[CFARUtils.scala 510:30]
  reg [31:0] _RAND_686;
  wire  cfar_cfar_cfarCore_leadWindow__T; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_1; // @[CFARUtils.scala 511:45]
  wire  cfar_cfar_cfarCore_leadWindow_en; // @[CFARUtils.scala 511:36]
  reg  cfar_cfar_cfarCore_leadWindow_validPrev; // @[CFARUtils.scala 514:26]
  reg [31:0] _RAND_687;
  wire [5:0] cfar_cfar_cfarCore_leadWindow__T_3; // @[CFARUtils.scala 515:21]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__GEN_140; // @[CFARUtils.scala 515:27]
  wire  cfar_cfar_cfarCore_leadWindow__T_4; // @[CFARUtils.scala 515:27]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__GEN_141; // @[CFARUtils.scala 516:28]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__T_6; // @[CFARUtils.scala 516:28]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__T_8; // @[CFARUtils.scala 516:39]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__T_10; // @[CFARUtils.scala 518:27]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__T_12; // @[CFARUtils.scala 518:41]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__T_14; // @[CFARUtils.scala 518:47]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__GEN_0; // @[CFARUtils.scala 515:40]
  wire [6:0] cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 528:34]
  wire  cfar_cfar_cfarCore_leadWindow__T_17; // @[CFARUtils.scala 528:21]
  wire  cfar_cfar_cfarCore_leadWindow__T_19; // @[CFARUtils.scala 528:40]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_1; // @[CFARUtils.scala 528:57]
  wire  cfar_cfar_cfarCore_leadWindow_fireLastIn; // @[CFARUtils.scala 531:30]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_2; // @[CFARUtils.scala 533:21]
  wire  cfar_cfar_cfarCore_leadWindow__T_21; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_22; // @[CFARUtils.scala 330:18]
  wire  cfar_cfar_cfarCore_leadWindow__T_24; // @[CFARUtils.scala 330:11]
  wire  cfar_cfar_cfarCore_leadWindow__T_25; // @[CFARUtils.scala 330:11]
  wire  cfar_cfar_cfarCore_leadWindow__T_33; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_37; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_41; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_45; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_49; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_53; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_57; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_61; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_65; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_69; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_73; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_77; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_81; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_85; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_89; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_93; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_97; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_101; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_105; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_109; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_113; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_117; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_121; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_125; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_129; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_133; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_137; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_141; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_145; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_149; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_153; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_157; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_161; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_165; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_169; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_173; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_177; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_181; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_185; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_189; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_193; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_197; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_201; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_205; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_209; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_213; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_217; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_221; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_225; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_229; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_233; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_237; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_241; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_245; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_249; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_253; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_257; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_261; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_265; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_269; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_273; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_277; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_281; // @[CFARUtils.scala 335:78]
  wire  cfar_cfar_cfarCore_leadWindow__T_284; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_285; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_286; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_287; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_288; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_289; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_290; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_291; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_292; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_293; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_294; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_295; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_296; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_297; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_298; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_299; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_300; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_301; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_302; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_303; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_304; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_305; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_306; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_307; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_308; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_309; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_310; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_311; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_312; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_313; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_314; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_315; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_316; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_317; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_318; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_319; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_320; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_321; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_322; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_323; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_324; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_325; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_326; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_327; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_328; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_329; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_330; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_331; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_332; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_333; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_334; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_335; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_336; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_337; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_338; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_339; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_340; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_341; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_342; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_343; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_344; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_345; // @[CFARUtils.scala 319:37]
  wire  cfar_cfar_cfarCore_leadWindow__T_346; // @[CFARUtils.scala 319:37]
  reg  cfar_cfar_cfarCore_leadWindow__T_348; // @[Reg.scala 27:20]
  reg [31:0] _RAND_688;
  reg  cfar_cfar_cfarCore_leadWindow__T_349; // @[Reg.scala 27:20]
  reg [31:0] _RAND_689;
  reg  cfar_cfar_cfarCore_leadWindow__T_350; // @[Reg.scala 27:20]
  reg [31:0] _RAND_690;
  reg  cfar_cfar_cfarCore_leadWindow__T_351; // @[Reg.scala 27:20]
  reg [31:0] _RAND_691;
  reg  cfar_cfar_cfarCore_leadWindow__T_352; // @[Reg.scala 27:20]
  reg [31:0] _RAND_692;
  reg  cfar_cfar_cfarCore_leadWindow__T_353; // @[Reg.scala 27:20]
  reg [31:0] _RAND_693;
  reg  cfar_cfar_cfarCore_leadWindow__T_354; // @[Reg.scala 27:20]
  reg [31:0] _RAND_694;
  reg  cfar_cfar_cfarCore_leadWindow__T_355; // @[Reg.scala 27:20]
  reg [31:0] _RAND_695;
  reg  cfar_cfar_cfarCore_leadWindow__T_356; // @[Reg.scala 27:20]
  reg [31:0] _RAND_696;
  reg  cfar_cfar_cfarCore_leadWindow__T_357; // @[Reg.scala 27:20]
  reg [31:0] _RAND_697;
  reg  cfar_cfar_cfarCore_leadWindow__T_358; // @[Reg.scala 27:20]
  reg [31:0] _RAND_698;
  reg  cfar_cfar_cfarCore_leadWindow__T_359; // @[Reg.scala 27:20]
  reg [31:0] _RAND_699;
  reg  cfar_cfar_cfarCore_leadWindow__T_360; // @[Reg.scala 27:20]
  reg [31:0] _RAND_700;
  reg  cfar_cfar_cfarCore_leadWindow__T_361; // @[Reg.scala 27:20]
  reg [31:0] _RAND_701;
  reg  cfar_cfar_cfarCore_leadWindow__T_362; // @[Reg.scala 27:20]
  reg [31:0] _RAND_702;
  reg  cfar_cfar_cfarCore_leadWindow__T_363; // @[Reg.scala 27:20]
  reg [31:0] _RAND_703;
  reg  cfar_cfar_cfarCore_leadWindow__T_364; // @[Reg.scala 27:20]
  reg [31:0] _RAND_704;
  reg  cfar_cfar_cfarCore_leadWindow__T_365; // @[Reg.scala 27:20]
  reg [31:0] _RAND_705;
  reg  cfar_cfar_cfarCore_leadWindow__T_366; // @[Reg.scala 27:20]
  reg [31:0] _RAND_706;
  reg  cfar_cfar_cfarCore_leadWindow__T_367; // @[Reg.scala 27:20]
  reg [31:0] _RAND_707;
  reg  cfar_cfar_cfarCore_leadWindow__T_368; // @[Reg.scala 27:20]
  reg [31:0] _RAND_708;
  reg  cfar_cfar_cfarCore_leadWindow__T_369; // @[Reg.scala 27:20]
  reg [31:0] _RAND_709;
  reg  cfar_cfar_cfarCore_leadWindow__T_370; // @[Reg.scala 27:20]
  reg [31:0] _RAND_710;
  reg  cfar_cfar_cfarCore_leadWindow__T_371; // @[Reg.scala 27:20]
  reg [31:0] _RAND_711;
  reg  cfar_cfar_cfarCore_leadWindow__T_372; // @[Reg.scala 27:20]
  reg [31:0] _RAND_712;
  reg  cfar_cfar_cfarCore_leadWindow__T_373; // @[Reg.scala 27:20]
  reg [31:0] _RAND_713;
  reg  cfar_cfar_cfarCore_leadWindow__T_374; // @[Reg.scala 27:20]
  reg [31:0] _RAND_714;
  reg  cfar_cfar_cfarCore_leadWindow__T_375; // @[Reg.scala 27:20]
  reg [31:0] _RAND_715;
  reg  cfar_cfar_cfarCore_leadWindow__T_376; // @[Reg.scala 27:20]
  reg [31:0] _RAND_716;
  reg  cfar_cfar_cfarCore_leadWindow__T_377; // @[Reg.scala 27:20]
  reg [31:0] _RAND_717;
  reg  cfar_cfar_cfarCore_leadWindow__T_378; // @[Reg.scala 27:20]
  reg [31:0] _RAND_718;
  reg  cfar_cfar_cfarCore_leadWindow__T_379; // @[Reg.scala 27:20]
  reg [31:0] _RAND_719;
  reg  cfar_cfar_cfarCore_leadWindow__T_380; // @[Reg.scala 27:20]
  reg [31:0] _RAND_720;
  reg  cfar_cfar_cfarCore_leadWindow__T_381; // @[Reg.scala 27:20]
  reg [31:0] _RAND_721;
  reg  cfar_cfar_cfarCore_leadWindow__T_382; // @[Reg.scala 27:20]
  reg [31:0] _RAND_722;
  reg  cfar_cfar_cfarCore_leadWindow__T_383; // @[Reg.scala 27:20]
  reg [31:0] _RAND_723;
  reg  cfar_cfar_cfarCore_leadWindow__T_384; // @[Reg.scala 27:20]
  reg [31:0] _RAND_724;
  reg  cfar_cfar_cfarCore_leadWindow__T_385; // @[Reg.scala 27:20]
  reg [31:0] _RAND_725;
  reg  cfar_cfar_cfarCore_leadWindow__T_386; // @[Reg.scala 27:20]
  reg [31:0] _RAND_726;
  reg  cfar_cfar_cfarCore_leadWindow__T_387; // @[Reg.scala 27:20]
  reg [31:0] _RAND_727;
  reg  cfar_cfar_cfarCore_leadWindow__T_388; // @[Reg.scala 27:20]
  reg [31:0] _RAND_728;
  reg  cfar_cfar_cfarCore_leadWindow__T_389; // @[Reg.scala 27:20]
  reg [31:0] _RAND_729;
  reg  cfar_cfar_cfarCore_leadWindow__T_390; // @[Reg.scala 27:20]
  reg [31:0] _RAND_730;
  reg  cfar_cfar_cfarCore_leadWindow__T_391; // @[Reg.scala 27:20]
  reg [31:0] _RAND_731;
  reg  cfar_cfar_cfarCore_leadWindow__T_392; // @[Reg.scala 27:20]
  reg [31:0] _RAND_732;
  reg  cfar_cfar_cfarCore_leadWindow__T_393; // @[Reg.scala 27:20]
  reg [31:0] _RAND_733;
  reg  cfar_cfar_cfarCore_leadWindow__T_394; // @[Reg.scala 27:20]
  reg [31:0] _RAND_734;
  reg  cfar_cfar_cfarCore_leadWindow__T_395; // @[Reg.scala 27:20]
  reg [31:0] _RAND_735;
  reg  cfar_cfar_cfarCore_leadWindow__T_396; // @[Reg.scala 27:20]
  reg [31:0] _RAND_736;
  reg  cfar_cfar_cfarCore_leadWindow__T_397; // @[Reg.scala 27:20]
  reg [31:0] _RAND_737;
  reg  cfar_cfar_cfarCore_leadWindow__T_398; // @[Reg.scala 27:20]
  reg [31:0] _RAND_738;
  reg  cfar_cfar_cfarCore_leadWindow__T_399; // @[Reg.scala 27:20]
  reg [31:0] _RAND_739;
  reg  cfar_cfar_cfarCore_leadWindow__T_400; // @[Reg.scala 27:20]
  reg [31:0] _RAND_740;
  reg  cfar_cfar_cfarCore_leadWindow__T_401; // @[Reg.scala 27:20]
  reg [31:0] _RAND_741;
  reg  cfar_cfar_cfarCore_leadWindow__T_402; // @[Reg.scala 27:20]
  reg [31:0] _RAND_742;
  reg  cfar_cfar_cfarCore_leadWindow__T_403; // @[Reg.scala 27:20]
  reg [31:0] _RAND_743;
  reg  cfar_cfar_cfarCore_leadWindow__T_404; // @[Reg.scala 27:20]
  reg [31:0] _RAND_744;
  reg  cfar_cfar_cfarCore_leadWindow__T_405; // @[Reg.scala 27:20]
  reg [31:0] _RAND_745;
  reg  cfar_cfar_cfarCore_leadWindow__T_406; // @[Reg.scala 27:20]
  reg [31:0] _RAND_746;
  reg  cfar_cfar_cfarCore_leadWindow__T_407; // @[Reg.scala 27:20]
  reg [31:0] _RAND_747;
  reg  cfar_cfar_cfarCore_leadWindow__T_408; // @[Reg.scala 27:20]
  reg [31:0] _RAND_748;
  reg  cfar_cfar_cfarCore_leadWindow__T_409; // @[Reg.scala 27:20]
  reg [31:0] _RAND_749;
  reg  cfar_cfar_cfarCore_leadWindow__T_410; // @[Reg.scala 27:20]
  reg [31:0] _RAND_750;
  reg  cfar_cfar_cfarCore_leadWindow__T_411; // @[Reg.scala 27:20]
  reg [31:0] _RAND_751;
  wire [5:0] cfar_cfar_cfarCore_leadWindow__T_414;
  wire  cfar_cfar_cfarCore_leadWindow__GEN_68; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_69; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_70; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_71; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_72; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_73; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_74; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_75; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_76; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_77; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_78; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_79; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_80; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_81; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_82; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_83; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_84; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_85; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_86; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_87; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_88; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_89; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_90; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_91; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_92; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_93; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_94; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_95; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_96; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_97; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_98; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_99; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_100; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_101; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_102; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_103; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_104; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_105; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_106; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_107; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_108; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_109; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_110; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_111; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_112; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_113; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_114; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_115; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_116; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_117; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_118; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_119; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_120; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_121; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_122; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_123; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_124; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_125; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_126; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_127; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_128; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_129; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__GEN_130; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow_resetAll; // @[CFARUtils.scala 537:26]
  wire  cfar_cfar_cfarCore_leadWindow__T_416; // @[CFARUtils.scala 544:15]
  wire  cfar_cfar_cfarCore_leadWindow__T_417; // @[CFARUtils.scala 544:12]
  wire  cfar_cfar_cfarCore_leadWindow__T_419; // @[CFARUtils.scala 546:36]
  reg [15:0] cfar_cfar_cfarCore_leadWindow__T_426; // @[CFARUtils.scala 551:37]
  reg [31:0] _RAND_752;
  wire  cfar_cfar_cfarCore_leadWindow__T_430; // @[CFARUtils.scala 554:31]
  wire  cfar_cfar_cfarCore_leadWindow__T_431; // @[CFARUtils.scala 554:42]
  wire  cfar_cfar_cfarCore_leadWindow__T_433; // @[CFARUtils.scala 555:36]
  wire  cfar_cfar_cfarCore_leadWindow__T_437; // @[CFARUtils.scala 568:33]
  wire  cfar_cfar_cfarCore_leadWindow__T_438; // @[CFARUtils.scala 568:57]
  wire [5:0] cfar_cfar_cfarCore_leadWindow_readIdx; // @[CFARUtils.scala 506:27 CFARUtils.scala 516:13 CFARUtils.scala 518:13]
  wire  cfar_cfar_cfarCore_Queue_clock;
  wire  cfar_cfar_cfarCore_Queue_reset;
  wire  cfar_cfar_cfarCore_Queue_io_enq_ready;
  wire  cfar_cfar_cfarCore_Queue_io_enq_valid;
  wire  cfar_cfar_cfarCore_Queue_io_enq_bits_peak;
  wire [15:0] cfar_cfar_cfarCore_Queue_io_enq_bits_cut;
  wire [15:0] cfar_cfar_cfarCore_Queue_io_enq_bits_threshold;
  wire  cfar_cfar_cfarCore_Queue_io_deq_ready;
  wire  cfar_cfar_cfarCore_Queue_io_deq_valid;
  wire  cfar_cfar_cfarCore_Queue_io_deq_bits_peak;
  wire [15:0] cfar_cfar_cfarCore_Queue_io_deq_bits_cut;
  wire [15:0] cfar_cfar_cfarCore_Queue_io_deq_bits_threshold;
  reg  cfar_cfar_cfarCore_Queue__T_peak [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_753;
  wire  cfar_cfar_cfarCore_Queue__T_peak__T_18_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_peak__T_18_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_peak__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_peak__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_peak__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_peak__T_10_en; // @[Decoupled.scala 209:24]
  reg [15:0] cfar_cfar_cfarCore_Queue__T_cut [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_754;
  wire [15:0] cfar_cfar_cfarCore_Queue__T_cut__T_18_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_cut__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] cfar_cfar_cfarCore_Queue__T_cut__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_cut__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_cut__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_cut__T_10_en; // @[Decoupled.scala 209:24]
  reg [15:0] cfar_cfar_cfarCore_Queue__T_threshold [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_755;
  wire [15:0] cfar_cfar_cfarCore_Queue__T_threshold__T_18_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_threshold__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] cfar_cfar_cfarCore_Queue__T_threshold__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_threshold__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_threshold__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue__T_threshold__T_10_en; // @[Decoupled.scala 209:24]
  reg  cfar_cfar_cfarCore_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_756;
  reg  cfar_cfar_cfarCore_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_757;
  reg  cfar_cfar_cfarCore_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_758;
  wire  cfar_cfar_cfarCore_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  cfar_cfar_cfarCore_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  cfar_cfar_cfarCore_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  cfar_cfar_cfarCore_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  cfar_cfar_cfarCore_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_Queue__T_12; // @[Counter.scala 39:22]
  wire  cfar_cfar_cfarCore_Queue__GEN_11; // @[Decoupled.scala 240:27]
  wire  cfar_cfar_cfarCore_Queue__GEN_16; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_Queue__T_14; // @[Counter.scala 39:22]
  wire  cfar_cfar_cfarCore_Queue__GEN_15; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_Queue__T_15; // @[Decoupled.scala 227:16]
  wire  cfar_cfar_cfarCore_Queue__T_16; // @[Decoupled.scala 231:19]
  wire  cfar_cfar_cfarCore_Queue_2_clock;
  wire  cfar_cfar_cfarCore_Queue_2_reset;
  wire  cfar_cfar_cfarCore_Queue_2_io_enq_ready;
  wire  cfar_cfar_cfarCore_Queue_2_io_enq_valid;
  wire  cfar_cfar_cfarCore_Queue_2_io_enq_bits;
  wire  cfar_cfar_cfarCore_Queue_2_io_deq_ready;
  wire  cfar_cfar_cfarCore_Queue_2_io_deq_valid;
  wire  cfar_cfar_cfarCore_Queue_2_io_deq_bits;
  reg  cfar_cfar_cfarCore_Queue_2__T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_759;
  wire  cfar_cfar_cfarCore_Queue_2__T__T_18_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue_2__T__T_18_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue_2__T__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue_2__T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue_2__T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_cfar_cfarCore_Queue_2__T__T_10_en; // @[Decoupled.scala 209:24]
  reg  cfar_cfar_cfarCore_Queue_2_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_760;
  reg  cfar_cfar_cfarCore_Queue_2_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_761;
  reg  cfar_cfar_cfarCore_Queue_2__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_762;
  wire  cfar_cfar_cfarCore_Queue_2__T_2; // @[Decoupled.scala 214:41]
  wire  cfar_cfar_cfarCore_Queue_2__T_3; // @[Decoupled.scala 215:36]
  wire  cfar_cfar_cfarCore_Queue_2__T_4; // @[Decoupled.scala 215:33]
  wire  cfar_cfar_cfarCore_Queue_2__T_5; // @[Decoupled.scala 216:32]
  wire  cfar_cfar_cfarCore_Queue_2__T_6; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_Queue_2__T_8; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore_Queue_2__T_12; // @[Counter.scala 39:22]
  wire  cfar_cfar_cfarCore_Queue_2__GEN_9; // @[Decoupled.scala 240:27]
  wire  cfar_cfar_cfarCore_Queue_2__GEN_12; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_Queue_2__T_14; // @[Counter.scala 39:22]
  wire  cfar_cfar_cfarCore_Queue_2__GEN_11; // @[Decoupled.scala 237:18]
  wire  cfar_cfar_cfarCore_Queue_2__T_15; // @[Decoupled.scala 227:16]
  wire  cfar_cfar_cfarCore_Queue_2__T_16; // @[Decoupled.scala 231:19]
  reg  cfar_cfar_cfarCore_lastCut; // @[CFARCoreWithMem.scala 20:24]
  reg [31:0] _RAND_763;
  reg  cfar_cfar_cfarCore_flushing; // @[CFARCoreWithMem.scala 21:25]
  reg [31:0] _RAND_764;
  reg [8:0] cfar_cfar_cfarCore_cntIn; // @[CFARCoreWithMem.scala 22:22]
  reg [31:0] _RAND_765;
  reg [8:0] cfar_cfar_cfarCore_cntOut; // @[CFARCoreWithMem.scala 23:23]
  reg [31:0] _RAND_766;
  reg  cfar_cfar_cfarCore_initialInDone; // @[CFARCoreWithMem.scala 24:30]
  reg [31:0] _RAND_767;
  wire [6:0] cfar_cfar_cfarCore__GEN_41; // @[CFARCoreWithMem.scala 32:32]
  wire [7:0] cfar_cfar_cfarCore__T; // @[CFARCoreWithMem.scala 32:32]
  wire [8:0] cfar_cfar_cfarCore_latency; // @[CFARCoreWithMem.scala 32:49]
  wire [8:0] cfar_cfar_cfarCore__T_1; // @[CFARCoreWithMem.scala 33:26]
  wire [5:0] cfar_cfar_cfarCore__T_2; // @[CFARCoreWithMem.scala 33:49]
  wire [8:0] cfar_cfar_cfarCore__GEN_42; // @[CFARCoreWithMem.scala 33:43]
  wire [8:0] cfar_cfar_cfarCore__T_4; // @[CFARCoreWithMem.scala 33:43]
  wire [8:0] cfar_cfar_cfarCore__T_6; // @[CFARCoreWithMem.scala 33:65]
  wire [9:0] cfar_cfar_cfarCore__GEN_43; // @[CFARCoreWithMem.scala 33:20]
  wire  cfar_cfar_cfarCore__T_7; // @[CFARCoreWithMem.scala 33:20]
  wire  cfar_cfar_cfarCore__T_9; // @[CFARCoreWithMem.scala 33:9]
  wire  cfar_cfar_cfarCore__T_10; // @[CFARCoreWithMem.scala 33:9]
  wire  cfar_cfar_cfarCore__T_11; // @[CFARCoreWithMem.scala 34:24]
  wire  cfar_cfar_cfarCore__T_13; // @[CFARCoreWithMem.scala 34:9]
  wire  cfar_cfar_cfarCore__T_14; // @[CFARCoreWithMem.scala 34:9]
  reg [19:0] cfar_cfar_cfarCore_sumlagg; // @[CFARCoreWithMem.scala 37:24]
  reg [31:0] _RAND_768;
  reg [19:0] cfar_cfar_cfarCore_sumlead; // @[CFARCoreWithMem.scala 38:24]
  reg [31:0] _RAND_769;
  reg  cfar_cfar_cfarCore_lastOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_770;
  wire  cfar_cfar_cfarCore__T_21; // @[Decoupled.scala 40:37]
  wire [8:0] cfar_cfar_cfarCore__T_23; // @[CFARCoreWithMem.scala 75:20]
  wire [8:0] cfar_cfar_cfarCore__T_25; // @[CFARCoreWithMem.scala 77:28]
  wire  cfar_cfar_cfarCore__T_26; // @[CFARCoreWithMem.scala 77:15]
  wire  cfar_cfar_cfarCore__T_28; // @[CFARCoreWithMem.scala 77:35]
  wire  cfar_cfar_cfarCore__GEN_2; // @[CFARCoreWithMem.scala 77:52]
  wire  cfar_cfar_cfarCore__T_29; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore__T_30; // @[CFARCoreWithMem.scala 81:20]
  wire [8:0] cfar_cfar_cfarCore__T_33; // @[CFARCoreWithMem.scala 85:22]
  wire [9:0] cfar_cfar_cfarCore__T_35; // @[CFARCoreWithMem.scala 87:31]
  wire [9:0] cfar_cfar_cfarCore__GEN_44; // @[CFARCoreWithMem.scala 87:16]
  wire  cfar_cfar_cfarCore__T_36; // @[CFARCoreWithMem.scala 87:16]
  wire  cfar_cfar_cfarCore__T_38; // @[CFARCoreWithMem.scala 87:38]
  wire  cfar_cfar_cfarCore__T_41; // @[CFARCoreWithMem.scala 87:55]
  wire  cfar_cfar_cfarCore__T_42; // @[CFARCoreWithMem.scala 93:19]
  wire  cfar_cfar_cfarCore__GEN_6; // @[CFARCoreWithMem.scala 93:35]
  reg  cfar_cfar_cfarCore_flushingDelayed; // @[CFARUtils.scala 286:20]
  reg [31:0] _RAND_771;
  wire  cfar_cfar_cfarCore__GEN_9; // @[CFARCoreWithMem.scala 101:21]
  wire  cfar_cfar_cfarCore__T_43; // @[CFARCoreWithMem.scala 106:32]
  wire  cfar_cfar_cfarCore__T_47; // @[Decoupled.scala 40:37]
  wire [19:0] cfar_cfar_cfarCore__GEN_45; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] cfar_cfar_cfarCore__T_50; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] cfar_cfar_cfarCore__GEN_46; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] cfar_cfar_cfarCore__T_53; // @[FixedPointTypeClass.scala 30:68]
  wire  cfar_cfar_cfarCore__T_59; // @[Decoupled.scala 40:37]
  wire  cfar_cfar_cfarCore__T_60; // @[Decoupled.scala 40:37]
  wire [19:0] cfar_cfar_cfarCore__GEN_48; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] cfar_cfar_cfarCore__T_63; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] cfar_cfar_cfarCore__GEN_49; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] cfar_cfar_cfarCore__T_66; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] cfar_cfar_cfarCore_leftThr; // @[FixedPointTypeClass.scala 118:51]
  wire [19:0] cfar_cfar_cfarCore_rightThr; // @[FixedPointTypeClass.scala 118:51]
  wire  cfar_cfar_cfarCore__T_70; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] cfar_cfar_cfarCore_greatestOf; // @[CFARCoreWithMem.scala 143:23]
  wire  cfar_cfar_cfarCore__T_71; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] cfar_cfar_cfarCore_smallestOf; // @[CFARCoreWithMem.scala 144:23]
  wire [19:0] cfar_cfar_cfarCore__T_74; // @[FixedPointTypeClass.scala 20:58]
  wire [18:0] cfar_cfar_cfarCore__T_75; // @[FixedPointTypeClass.scala 117:50]
  wire  cfar_cfar_cfarCore__T_78; // @[Mux.scala 68:19]
  wire [19:0] cfar_cfar_cfarCore__T_79; // @[Mux.scala 68:16]
  wire  cfar_cfar_cfarCore__T_80; // @[Mux.scala 68:19]
  wire [19:0] cfar_cfar_cfarCore_thrByModes; // @[Mux.scala 68:16]
  reg  cfar_cfar_cfarCore_enableRightThr; // @[CFARCoreWithMem.scala 151:31]
  reg [31:0] _RAND_772;
  wire  cfar_cfar_cfarCore__T_81; // @[CFARCoreWithMem.scala 152:9]
  wire  cfar_cfar_cfarCore__T_83; // @[CFARCoreWithMem.scala 152:34]
  wire  cfar_cfar_cfarCore__GEN_21; // @[CFARCoreWithMem.scala 152:63]
  wire  cfar_cfar_cfarCore__T_84; // @[CFARCoreWithMem.scala 172:33]
  wire  cfar_cfar_cfarCore__T_86; // @[CFARCoreWithMem.scala 172:56]
  wire  cfar_cfar_cfarCore__T_90; // @[CFARCoreWithMem.scala 174:57]
  wire [19:0] cfar_cfar_cfarCore__T_91; // @[CFARCoreWithMem.scala 177:36]
  wire [19:0] cfar_cfar_cfarCore__T_92; // @[CFARCoreWithMem.scala 174:34]
  wire [19:0] cfar_cfar_cfarCore_thrWithoutScaling; // @[CFARCoreWithMem.scala 172:32]
  wire [19:0] cfar_cfar_cfarCore__GEN_51; // @[FixedPointTypeClass.scala 211:35]
  reg [35:0] cfar_cfar_cfarCore__T_94; // @[Reg.scala 15:16]
  reg [63:0] _RAND_773;
  wire [22:0] cfar_cfar_cfarCore_threshold; // @[FixedPointTypeClass.scala 153:43]
  reg [15:0] cfar_cfar_cfarCore_cutDelayed; // @[Reg.scala 15:16]
  reg [31:0] _RAND_774;
  wire [3:0] cfar_cfar_cfarCore__T_96; // @[CFARCoreWithMem.scala 197:74]
  wire [2:0] cfar_cfar_cfarCore__T_97;
  reg [15:0] cfar_cfar_cfarCore_leftNeighb; // @[Reg.scala 15:16]
  reg [31:0] _RAND_775;
  wire [15:0] cfar_cfar_cfarCore__GEN_25; // @[Reg.scala 16:23]
  reg [15:0] cfar_cfar_cfarCore_rightNeighb; // @[Reg.scala 15:16]
  reg [31:0] _RAND_776;
  wire  cfar_cfar_cfarCore__T_98; // @[FixedPointTypeClass.scala 55:59]
  wire  cfar_cfar_cfarCore__T_99; // @[FixedPointTypeClass.scala 55:59]
  wire  cfar_cfar_cfarCore_isLocalMax; // @[CFARCoreWithMem.scala 199:44]
  wire [16:0] cfar_cfar_cfarCore__GEN_52; // @[FixedPointTypeClass.scala 55:59]
  wire [22:0] cfar_cfar_cfarCore__GEN_53; // @[FixedPointTypeClass.scala 55:59]
  wire  cfar_cfar_cfarCore_isPeak; // @[FixedPointTypeClass.scala 55:59]
  wire  cfar_cfar_cfarCore__T_100; // @[CFARCoreWithMem.scala 216:20]
  wire  cfar_cfar_cfarCore__T_101; // @[CFARCoreWithMem.scala 216:54]
  wire  cfar_cfar_cfarCore__T_102; // @[CFARCoreWithMem.scala 216:51]
  reg  cfar_cfar_cfarCore__T_106; // @[Reg.scala 15:16]
  reg [31:0] _RAND_777;
  reg  cfar_cfar_cfarCore__T_107; // @[Reg.scala 15:16]
  reg [31:0] _RAND_778;
  wire  cfar_cfar_cfarCore__T_108; // @[CFARCoreWithMem.scala 218:123]
  wire  cfar_cfar_cfarCore__T_110; // @[CFARCoreWithMem.scala 223:63]
  reg  cfar_cfar_cfarCore__T_120; // @[Reg.scala 15:16]
  reg [31:0] _RAND_779;
  reg  cfar_cfar_cfarCore__T_121; // @[Reg.scala 15:16]
  reg [31:0] _RAND_780;
  wire  cfar_cfar_cfarCore__T_122; // @[CFARCoreWithMem.scala 231:123]
  wire [21:0] cfar_cfar_cfarCore__GEN_55; // @[CFARCoreWithMem.scala 222:37]
  wire  cfar_Queue_clock;
  wire  cfar_Queue_reset;
  wire  cfar_Queue_io_enq_ready;
  wire  cfar_Queue_io_enq_valid;
  wire  cfar_Queue_io_enq_bits_read;
  wire [31:0] cfar_Queue_io_enq_bits_data;
  wire  cfar_Queue_io_enq_bits_extra;
  wire  cfar_Queue_io_deq_ready;
  wire  cfar_Queue_io_deq_valid;
  wire  cfar_Queue_io_deq_bits_read;
  wire [31:0] cfar_Queue_io_deq_bits_data;
  wire  cfar_Queue_io_deq_bits_extra;
  reg  cfar_Queue__T_read [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_781;
  wire  cfar_Queue__T_read__T_18_data; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_read__T_18_addr; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_read__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_read__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_read__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_read__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] cfar_Queue__T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_782;
  wire [31:0] cfar_Queue__T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] cfar_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  cfar_Queue__T_extra [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_783;
  wire  cfar_Queue__T_extra__T_18_data; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_extra__T_18_addr; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_extra__T_10_data; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_extra__T_10_addr; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_extra__T_10_mask; // @[Decoupled.scala 209:24]
  wire  cfar_Queue__T_extra__T_10_en; // @[Decoupled.scala 209:24]
  reg  cfar_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_784;
  reg  cfar_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_785;
  reg  cfar_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_786;
  wire  cfar_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  cfar_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  cfar_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  cfar_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  cfar_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  cfar_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  cfar_Queue__T_12; // @[Counter.scala 39:22]
  wire  cfar_Queue__T_14; // @[Counter.scala 39:22]
  wire  cfar_Queue__T_15; // @[Decoupled.scala 227:16]
  reg [9:0] cfar_fftWin; // @[CFARDspBlock.scala 72:25]
  reg [31:0] _RAND_787;
  reg [15:0] cfar_thresholdScaler; // @[CFARDspBlock.scala 73:34]
  reg [31:0] _RAND_788;
  reg  cfar_peakGrouping; // @[CFARDspBlock.scala 74:31]
  reg [31:0] _RAND_789;
  reg [1:0] cfar_cfarMode; // @[CFARDspBlock.scala 75:27]
  reg [31:0] _RAND_790;
  reg [6:0] cfar_windowCells; // @[CFARDspBlock.scala 76:30]
  reg [31:0] _RAND_791;
  reg [3:0] cfar_guardCells; // @[CFARDspBlock.scala 77:29]
  reg [31:0] _RAND_792;
  reg [2:0] cfar__T_6; // @[CFARDspBlock.scala 111:27]
  reg [31:0] _RAND_793;
  wire [41:0] cfar__T_11; // @[Cat.scala 29:58]
  wire  cfar__T_13; // @[RegisterRouter.scala 40:39]
  wire  cfar__T_14; // @[RegisterRouter.scala 40:26]
  wire  cfar__T_15; // @[RegisterRouter.scala 42:29]
  wire  cfar__T_58_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] cfar__T_22; // @[RegisterRouter.scala 48:19]
  wire [27:0] cfar__T_56; // @[RegisterRouter.scala 52:27]
  wire [5:0] cfar__T_12_bits_index; // @[RegisterRouter.scala 37:18 RegisterRouter.scala 52:19]
  wire  cfar__T_282; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_281; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_280; // @[RegisterRouter.scala 59:16]
  wire [2:0] cfar__T_287; // @[Cat.scala 29:58]
  wire [5:0] cfar__T_62; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_70; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_16; // @[RegisterRouter.scala 42:26]
  wire  cfar__T_24; // @[OneHot.scala 64:49]
  wire [1:0] cfar__T_25; // @[OneHot.scala 65:12]
  wire [1:0] cfar__T_27; // @[Misc.scala 200:81]
  wire  cfar__T_28; // @[Misc.scala 204:21]
  wire  cfar__T_29; // @[Misc.scala 207:26]
  wire  cfar__T_30; // @[Misc.scala 208:26]
  wire  cfar__T_31; // @[Misc.scala 209:20]
  wire  cfar__T_33; // @[Misc.scala 213:38]
  wire  cfar__T_34; // @[Misc.scala 213:29]
  wire  cfar__T_36; // @[Misc.scala 213:38]
  wire  cfar__T_37; // @[Misc.scala 213:29]
  wire  cfar__T_38; // @[Misc.scala 207:26]
  wire  cfar__T_39; // @[Misc.scala 208:26]
  wire  cfar__T_40; // @[Misc.scala 209:20]
  wire  cfar__T_41; // @[Misc.scala 212:27]
  wire  cfar__T_42; // @[Misc.scala 213:38]
  wire  cfar__T_43; // @[Misc.scala 213:29]
  wire  cfar__T_44; // @[Misc.scala 212:27]
  wire  cfar__T_45; // @[Misc.scala 213:38]
  wire  cfar__T_46; // @[Misc.scala 213:29]
  wire  cfar__T_47; // @[Misc.scala 212:27]
  wire  cfar__T_48; // @[Misc.scala 213:38]
  wire  cfar__T_49; // @[Misc.scala 213:29]
  wire  cfar__T_50; // @[Misc.scala 212:27]
  wire  cfar__T_51; // @[Misc.scala 213:38]
  wire  cfar__T_52; // @[Misc.scala 213:29]
  wire [3:0] cfar__T_55; // @[Cat.scala 29:58]
  wire [3:0] cfar__T_57; // @[RegisterRouter.scala 54:25]
  wire  cfar__T_81; // @[Bitwise.scala 26:51]
  wire  cfar__T_82; // @[Bitwise.scala 26:51]
  wire  cfar__T_83; // @[Bitwise.scala 26:51]
  wire  cfar__T_84; // @[Bitwise.scala 26:51]
  wire [7:0] cfar__T_86; // @[Bitwise.scala 72:12]
  wire [7:0] cfar__T_88; // @[Bitwise.scala 72:12]
  wire [7:0] cfar__T_90; // @[Bitwise.scala 72:12]
  wire [7:0] cfar__T_92; // @[Bitwise.scala 72:12]
  wire [31:0] cfar__T_95; // @[Cat.scala 29:58]
  wire [9:0] cfar__T_111; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_114; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_306; // @[RegisterRouter.scala 59:16]
  wire [7:0] cfar__T_288; // @[OneHot.scala 58:35]
  wire  cfar__T_289; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_353; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_355; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_356; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_121; // @[RegisterRouter.scala 59:16]
  wire [9:0] cfar__T_123; // @[RegisterRouter.scala 59:16]
  wire [3:0] cfar__T_134; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_137; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_294; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_380; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_381; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_144; // @[RegisterRouter.scala 59:16]
  wire [3:0] cfar__T_146; // @[RegisterRouter.scala 59:16]
  wire [15:0] cfar__T_157; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_160; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_290; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_360; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_361; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_167; // @[RegisterRouter.scala 59:16]
  wire [15:0] cfar__T_169; // @[RegisterRouter.scala 59:16]
  wire [2:0] cfar__T_180; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_183; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_295; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_385; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_386; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_190; // @[RegisterRouter.scala 59:16]
  wire [2:0] cfar__T_192; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_203; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_291; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_365; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_366; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_213; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_215; // @[RegisterRouter.scala 59:16]
  wire [1:0] cfar__T_226; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_229; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_292; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_370; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_371; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_236; // @[RegisterRouter.scala 59:16]
  wire [1:0] cfar__T_238; // @[RegisterRouter.scala 59:16]
  wire [6:0] cfar__T_249; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_252; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_293; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_375; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_376; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_259; // @[RegisterRouter.scala 59:16]
  wire [6:0] cfar__T_261; // @[RegisterRouter.scala 59:16]
  wire  cfar__GEN_40; // @[MuxLiteral.scala 48:10]
  wire  cfar__GEN_41; // @[MuxLiteral.scala 48:10]
  wire  cfar__GEN_42; // @[MuxLiteral.scala 48:10]
  wire  cfar__GEN_43; // @[MuxLiteral.scala 48:10]
  wire  cfar__GEN_44; // @[MuxLiteral.scala 48:10]
  wire  cfar__GEN_45; // @[MuxLiteral.scala 48:10]
  wire  cfar__GEN_55; // @[MuxLiteral.scala 48:10]
  wire  cfar__GEN_46; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__T_498_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] cfar__GEN_48; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__T_498_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] cfar__GEN_49; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__T_498_3; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] cfar__GEN_50; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__T_498_4; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] cfar__GEN_51; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__T_498_5; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] cfar__GEN_52; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__T_498_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] cfar__GEN_53; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__GEN_54; // @[MuxLiteral.scala 48:10]
  wire [15:0] cfar__T_500; // @[RegisterRouter.scala 59:16]
  wire  cfar__T_501_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  cfar__T_501_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  cfar__T_504; // @[RegisterRouter.scala 65:29]
  wire  widthAdapter_1_clock;
  wire  widthAdapter_1_reset;
  wire  widthAdapter_1_auto_in_ready;
  wire  widthAdapter_1_auto_in_valid;
  wire [47:0] widthAdapter_1_auto_in_bits_data;
  wire  widthAdapter_1_auto_in_bits_last;
  wire  widthAdapter_1_auto_out_ready;
  wire  widthAdapter_1_auto_out_valid;
  wire [15:0] widthAdapter_1_auto_out_bits_data;
  wire  widthAdapter_1_auto_out_bits_last;
  wire [15:0] widthAdapter_1__T; // @[AXI4StreamWidthAdapter.scala 154:10]
  wire [15:0] widthAdapter_1__T_1; // @[AXI4StreamWidthAdapter.scala 154:10]
  wire [15:0] widthAdapter_1__T_2; // @[AXI4StreamWidthAdapter.scala 154:10]
  reg [1:0] widthAdapter_1__T_4; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_794;
  wire  widthAdapter_1__T_5; // @[AXI4StreamWidthAdapter.scala 159:14]
  wire  widthAdapter_1__T_6; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] widthAdapter_1__T_7; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] widthAdapter_1__T_8; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] widthAdapter_1__GEN_0; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  widthAdapter_1_ir0; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] widthAdapter_1__T_10; // @[AXI4StreamWidthAdapter.scala 167:22]
  reg [31:0] _RAND_795;
  wire  widthAdapter_1__T_12; // @[AXI4StreamWidthAdapter.scala 168:38]
  wire [2:0] widthAdapter_1__T_13; // @[AXI4StreamWidthAdapter.scala 168:60]
  wire [2:0] widthAdapter_1__T_14; // @[AXI4StreamWidthAdapter.scala 168:33]
  wire [2:0] widthAdapter_1__GEN_1; // @[AXI4StreamWidthAdapter.scala 168:21]
  wire  widthAdapter_1_ir1; // @[AXI4StreamWidthAdapter.scala 170:60]
  reg [1:0] widthAdapter_1__T_19; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_796;
  wire  widthAdapter_1__T_21; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] widthAdapter_1__T_22; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] widthAdapter_1__T_23; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] widthAdapter_1__GEN_2; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  widthAdapter_1_ir2; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] widthAdapter_1__T_26; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_797;
  wire  widthAdapter_1__T_28; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] widthAdapter_1__T_29; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] widthAdapter_1__T_30; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] widthAdapter_1__GEN_3; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  widthAdapter_1_ir3; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] widthAdapter_1__T_33; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_798;
  wire  widthAdapter_1__T_35; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] widthAdapter_1__T_36; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] widthAdapter_1__T_37; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] widthAdapter_1__GEN_4; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  widthAdapter_1_ir4; // @[AXI4StreamWidthAdapter.scala 163:34]
  wire  widthAdapter_1__T_55; // @[AXI4StreamWidthAdapter.scala 46:16]
  wire  widthAdapter_1__T_57; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  widthAdapter_1__T_58; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  widthAdapter_1__T_59; // @[AXI4StreamWidthAdapter.scala 47:16]
  wire  widthAdapter_1__T_61; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  widthAdapter_1__T_62; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  widthAdapter_1__T_63; // @[AXI4StreamWidthAdapter.scala 48:16]
  wire  widthAdapter_1__T_65; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  widthAdapter_1__T_66; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  widthAdapter_1__T_67; // @[AXI4StreamWidthAdapter.scala 49:16]
  wire  widthAdapter_1__T_69; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire  widthAdapter_1__T_70; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire [15:0] widthAdapter_1__GEN_6; // @[AXI4StreamWidthAdapter.scala 54:19]
  wire  buffer_clock;
  wire  buffer_reset;
  wire  buffer_auto_in_ready;
  wire  buffer_auto_in_valid;
  wire [31:0] buffer_auto_in_bits_data;
  wire  buffer_auto_in_bits_last;
  wire  buffer_auto_out_ready;
  wire  buffer_auto_out_valid;
  wire [31:0] buffer_auto_out_bits_data;
  wire  buffer_auto_out_bits_last;
  wire  buffer_Queue_clock;
  wire  buffer_Queue_reset;
  wire  buffer_Queue_io_enq_ready;
  wire  buffer_Queue_io_enq_valid;
  wire [31:0] buffer_Queue_io_enq_bits_data;
  wire  buffer_Queue_io_enq_bits_last;
  wire  buffer_Queue_io_deq_ready;
  wire  buffer_Queue_io_deq_valid;
  wire [31:0] buffer_Queue_io_deq_bits_data;
  wire  buffer_Queue_io_deq_bits_last;
  reg [31:0] buffer_Queue__T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_799;
  wire [31:0] buffer_Queue__T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] buffer_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_Queue__T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_800;
  wire  buffer_Queue__T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_Queue__T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_801;
  reg  buffer_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_802;
  reg  buffer_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_803;
  wire  buffer_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  buffer_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  buffer_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  buffer_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  buffer_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  buffer_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  buffer_Queue__T_12; // @[Counter.scala 39:22]
  wire  buffer_Queue__T_14; // @[Counter.scala 39:22]
  wire  buffer_Queue__T_15; // @[Decoupled.scala 227:16]
  wire  buffer_1_clock;
  wire  buffer_1_reset;
  wire  buffer_1_auto_in_ready;
  wire  buffer_1_auto_in_valid;
  wire [15:0] buffer_1_auto_in_bits_data;
  wire  buffer_1_auto_in_bits_last;
  wire  buffer_1_auto_out_ready;
  wire  buffer_1_auto_out_valid;
  wire [15:0] buffer_1_auto_out_bits_data;
  wire  buffer_1_auto_out_bits_last;
  wire  buffer_1_Queue_clock;
  wire  buffer_1_Queue_reset;
  wire  buffer_1_Queue_io_enq_ready;
  wire  buffer_1_Queue_io_enq_valid;
  wire [15:0] buffer_1_Queue_io_enq_bits_data;
  wire  buffer_1_Queue_io_enq_bits_last;
  wire  buffer_1_Queue_io_deq_ready;
  wire  buffer_1_Queue_io_deq_valid;
  wire [15:0] buffer_1_Queue_io_deq_bits_data;
  wire  buffer_1_Queue_io_deq_bits_last;
  reg [15:0] buffer_1_Queue__T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_804;
  wire [15:0] buffer_1_Queue__T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] buffer_1_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_1_Queue__T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_805;
  wire  buffer_1_Queue__T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_1_Queue__T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_1_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_806;
  reg  buffer_1_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_807;
  reg  buffer_1_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_808;
  wire  buffer_1_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  buffer_1_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  buffer_1_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  buffer_1_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  buffer_1_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  buffer_1_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  buffer_1_Queue__T_12; // @[Counter.scala 39:22]
  wire  buffer_1_Queue__T_14; // @[Counter.scala 39:22]
  wire  buffer_1_Queue__T_15; // @[Decoupled.scala 227:16]
  wire  buffer_2_clock;
  wire  buffer_2_reset;
  wire  buffer_2_auto_in_ready;
  wire  buffer_2_auto_in_valid;
  wire [31:0] buffer_2_auto_in_bits_data;
  wire  buffer_2_auto_in_bits_last;
  wire  buffer_2_auto_out_ready;
  wire  buffer_2_auto_out_valid;
  wire [31:0] buffer_2_auto_out_bits_data;
  wire  buffer_2_auto_out_bits_last;
  wire  buffer_2_Queue_clock;
  wire  buffer_2_Queue_reset;
  wire  buffer_2_Queue_io_enq_ready;
  wire  buffer_2_Queue_io_enq_valid;
  wire [31:0] buffer_2_Queue_io_enq_bits_data;
  wire  buffer_2_Queue_io_enq_bits_last;
  wire  buffer_2_Queue_io_deq_ready;
  wire  buffer_2_Queue_io_deq_valid;
  wire [31:0] buffer_2_Queue_io_deq_bits_data;
  wire  buffer_2_Queue_io_deq_bits_last;
  reg [31:0] buffer_2_Queue__T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_809;
  wire [31:0] buffer_2_Queue__T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] buffer_2_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_2_Queue__T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_810;
  wire  buffer_2_Queue__T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_2_Queue__T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_2_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_811;
  reg  buffer_2_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_812;
  reg  buffer_2_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_813;
  wire  buffer_2_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  buffer_2_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  buffer_2_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  buffer_2_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  buffer_2_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  buffer_2_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  buffer_2_Queue__T_12; // @[Counter.scala 39:22]
  wire  buffer_2_Queue__T_14; // @[Counter.scala 39:22]
  wire  buffer_2_Queue__T_15; // @[Decoupled.scala 227:16]
  wire  buffer_3_clock;
  wire  buffer_3_reset;
  wire  buffer_3_auto_in_ready;
  wire  buffer_3_auto_in_valid;
  wire [47:0] buffer_3_auto_in_bits_data;
  wire  buffer_3_auto_in_bits_last;
  wire  buffer_3_auto_out_ready;
  wire  buffer_3_auto_out_valid;
  wire [47:0] buffer_3_auto_out_bits_data;
  wire  buffer_3_auto_out_bits_last;
  wire  buffer_3_Queue_clock;
  wire  buffer_3_Queue_reset;
  wire  buffer_3_Queue_io_enq_ready;
  wire  buffer_3_Queue_io_enq_valid;
  wire [47:0] buffer_3_Queue_io_enq_bits_data;
  wire  buffer_3_Queue_io_enq_bits_last;
  wire  buffer_3_Queue_io_deq_ready;
  wire  buffer_3_Queue_io_deq_valid;
  wire [47:0] buffer_3_Queue_io_deq_bits_data;
  wire  buffer_3_Queue_io_deq_bits_last;
  reg [47:0] buffer_3_Queue__T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [63:0] _RAND_814;
  wire [47:0] buffer_3_Queue__T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [47:0] buffer_3_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_3_Queue__T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_815;
  wire  buffer_3_Queue__T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  buffer_3_Queue__T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  buffer_3_Queue_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_816;
  reg  buffer_3_Queue_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_817;
  reg  buffer_3_Queue__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_818;
  wire  buffer_3_Queue__T_2; // @[Decoupled.scala 214:41]
  wire  buffer_3_Queue__T_3; // @[Decoupled.scala 215:36]
  wire  buffer_3_Queue__T_4; // @[Decoupled.scala 215:33]
  wire  buffer_3_Queue__T_5; // @[Decoupled.scala 216:32]
  wire  buffer_3_Queue__T_6; // @[Decoupled.scala 40:37]
  wire  buffer_3_Queue__T_8; // @[Decoupled.scala 40:37]
  wire  buffer_3_Queue__T_12; // @[Counter.scala 39:22]
  wire  buffer_3_Queue__T_14; // @[Counter.scala 39:22]
  wire  buffer_3_Queue__T_15; // @[Decoupled.scala 227:16]
  wire  bus_clock;
  wire  bus_reset;
  wire  bus_auto_in_aw_ready;
  wire  bus_auto_in_aw_valid;
  wire  bus_auto_in_aw_bits_id;
  wire [29:0] bus_auto_in_aw_bits_addr;
  wire  bus_auto_in_w_ready;
  wire  bus_auto_in_w_valid;
  wire [31:0] bus_auto_in_w_bits_data;
  wire [3:0] bus_auto_in_w_bits_strb;
  wire  bus_auto_in_w_bits_last;
  wire  bus_auto_in_b_ready;
  wire  bus_auto_in_b_valid;
  wire [1:0] bus_auto_in_b_bits_resp;
  wire  bus_auto_in_ar_ready;
  wire  bus_auto_in_ar_valid;
  wire  bus_auto_in_ar_bits_id;
  wire [29:0] bus_auto_in_ar_bits_addr;
  wire [2:0] bus_auto_in_ar_bits_size;
  wire  bus_auto_in_r_ready;
  wire  bus_auto_in_r_valid;
  wire [31:0] bus_auto_in_r_bits_data;
  wire [1:0] bus_auto_in_r_bits_resp;
  wire  bus_auto_in_r_bits_last;
  wire  bus_auto_out_2_aw_ready;
  wire  bus_auto_out_2_aw_valid;
  wire  bus_auto_out_2_aw_bits_id;
  wire [29:0] bus_auto_out_2_aw_bits_addr;
  wire  bus_auto_out_2_w_ready;
  wire  bus_auto_out_2_w_valid;
  wire [31:0] bus_auto_out_2_w_bits_data;
  wire [3:0] bus_auto_out_2_w_bits_strb;
  wire  bus_auto_out_2_b_ready;
  wire  bus_auto_out_2_b_valid;
  wire  bus_auto_out_2_b_bits_id;
  wire  bus_auto_out_2_ar_ready;
  wire  bus_auto_out_2_ar_valid;
  wire  bus_auto_out_2_ar_bits_id;
  wire [29:0] bus_auto_out_2_ar_bits_addr;
  wire [2:0] bus_auto_out_2_ar_bits_size;
  wire  bus_auto_out_2_r_ready;
  wire  bus_auto_out_2_r_valid;
  wire  bus_auto_out_2_r_bits_id;
  wire [31:0] bus_auto_out_2_r_bits_data;
  wire  bus_auto_out_1_aw_ready;
  wire  bus_auto_out_1_aw_valid;
  wire  bus_auto_out_1_aw_bits_id;
  wire [29:0] bus_auto_out_1_aw_bits_addr;
  wire  bus_auto_out_1_w_ready;
  wire  bus_auto_out_1_w_valid;
  wire [31:0] bus_auto_out_1_w_bits_data;
  wire [3:0] bus_auto_out_1_w_bits_strb;
  wire  bus_auto_out_1_b_ready;
  wire  bus_auto_out_1_b_valid;
  wire  bus_auto_out_1_b_bits_id;
  wire  bus_auto_out_1_ar_ready;
  wire  bus_auto_out_1_ar_valid;
  wire  bus_auto_out_1_ar_bits_id;
  wire [29:0] bus_auto_out_1_ar_bits_addr;
  wire [2:0] bus_auto_out_1_ar_bits_size;
  wire  bus_auto_out_1_r_ready;
  wire  bus_auto_out_1_r_valid;
  wire  bus_auto_out_1_r_bits_id;
  wire [31:0] bus_auto_out_1_r_bits_data;
  wire  bus_auto_out_0_aw_ready;
  wire  bus_auto_out_0_aw_valid;
  wire  bus_auto_out_0_aw_bits_id;
  wire [29:0] bus_auto_out_0_aw_bits_addr;
  wire  bus_auto_out_0_w_ready;
  wire  bus_auto_out_0_w_valid;
  wire  bus_auto_out_0_b_ready;
  wire  bus_auto_out_0_b_valid;
  wire  bus_auto_out_0_b_bits_id;
  wire  bus_auto_out_0_ar_ready;
  wire  bus_auto_out_0_ar_valid;
  wire  bus_auto_out_0_ar_bits_id;
  wire [29:0] bus_auto_out_0_ar_bits_addr;
  wire  bus_auto_out_0_r_ready;
  wire  bus_auto_out_0_r_valid;
  wire  bus_auto_out_0_r_bits_id;
  wire [31:0] bus_auto_out_0_r_bits_data;
  wire  bus_awIn_0_clock;
  wire  bus_awIn_0_reset;
  wire  bus_awIn_0_io_enq_ready;
  wire  bus_awIn_0_io_enq_valid;
  wire [2:0] bus_awIn_0_io_enq_bits;
  wire  bus_awIn_0_io_deq_ready;
  wire  bus_awIn_0_io_deq_valid;
  wire [2:0] bus_awIn_0_io_deq_bits;
  reg [2:0] bus_awIn_0__T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_819;
  wire [2:0] bus_awIn_0__T__T_18_data; // @[Decoupled.scala 209:24]
  wire  bus_awIn_0__T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [2:0] bus_awIn_0__T__T_10_data; // @[Decoupled.scala 209:24]
  wire  bus_awIn_0__T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  bus_awIn_0__T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  bus_awIn_0__T__T_10_en; // @[Decoupled.scala 209:24]
  reg  bus_awIn_0_value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_820;
  reg  bus_awIn_0_value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_821;
  reg  bus_awIn_0__T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_822;
  wire  bus_awIn_0__T_2; // @[Decoupled.scala 214:41]
  wire  bus_awIn_0__T_3; // @[Decoupled.scala 215:36]
  wire  bus_awIn_0__T_4; // @[Decoupled.scala 215:33]
  wire  bus_awIn_0__T_5; // @[Decoupled.scala 216:32]
  wire  bus_awIn_0__T_6; // @[Decoupled.scala 40:37]
  wire  bus_awIn_0__T_8; // @[Decoupled.scala 40:37]
  wire  bus_awIn_0__T_12; // @[Counter.scala 39:22]
  wire  bus_awIn_0__GEN_9; // @[Decoupled.scala 240:27]
  wire  bus_awIn_0__GEN_12; // @[Decoupled.scala 237:18]
  wire  bus_awIn_0__T_14; // @[Counter.scala 39:22]
  wire  bus_awIn_0__GEN_11; // @[Decoupled.scala 237:18]
  wire  bus_awIn_0__T_15; // @[Decoupled.scala 227:16]
  wire  bus_awIn_0__T_16; // @[Decoupled.scala 231:19]
  wire [30:0] bus__T_1; // @[Parameters.scala 137:49]
  wire [30:0] bus__T_3; // @[Parameters.scala 137:52]
  wire  bus_requestARIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] bus__T_5; // @[Parameters.scala 137:31]
  wire [30:0] bus__T_6; // @[Parameters.scala 137:49]
  wire [30:0] bus__T_8; // @[Parameters.scala 137:52]
  wire  bus_requestARIO_0_1; // @[Parameters.scala 137:67]
  wire [29:0] bus__T_10; // @[Parameters.scala 137:31]
  wire [30:0] bus__T_11; // @[Parameters.scala 137:49]
  wire [30:0] bus__T_13; // @[Parameters.scala 137:52]
  wire  bus_requestARIO_0_2; // @[Parameters.scala 137:67]
  wire [30:0] bus__T_16; // @[Parameters.scala 137:49]
  wire [30:0] bus__T_18; // @[Parameters.scala 137:52]
  wire  bus_requestAWIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] bus__T_20; // @[Parameters.scala 137:31]
  wire [30:0] bus__T_21; // @[Parameters.scala 137:49]
  wire [30:0] bus__T_23; // @[Parameters.scala 137:52]
  wire  bus_requestAWIO_0_1; // @[Parameters.scala 137:67]
  wire [29:0] bus__T_25; // @[Parameters.scala 137:31]
  wire [30:0] bus__T_26; // @[Parameters.scala 137:49]
  wire [30:0] bus__T_28; // @[Parameters.scala 137:52]
  wire  bus_requestAWIO_0_2; // @[Parameters.scala 137:67]
  wire  bus_requestROI_0_0; // @[Parameters.scala 47:9]
  wire  bus_requestROI_1_0; // @[Parameters.scala 47:9]
  wire  bus_requestROI_2_0; // @[Parameters.scala 47:9]
  wire  bus_requestBOI_0_0; // @[Parameters.scala 47:9]
  wire  bus_requestBOI_1_0; // @[Parameters.scala 47:9]
  wire  bus_requestBOI_2_0; // @[Parameters.scala 47:9]
  wire [1:0] bus__T_30; // @[Xbar.scala 64:75]
  wire [2:0] bus__T_31; // @[Xbar.scala 64:75]
  wire  bus_requestWIO_0_0; // @[Xbar.scala 65:73]
  wire  bus_requestWIO_0_1; // @[Xbar.scala 65:73]
  wire  bus_requestWIO_0_2; // @[Xbar.scala 65:73]
  wire [2:0] bus__T_39; // @[Xbar.scala 93:45]
  wire  bus__T_40; // @[OneHot.scala 30:18]
  wire [1:0] bus__T_41; // @[OneHot.scala 31:18]
  wire [1:0] bus__GEN_22; // @[OneHot.scala 32:28]
  wire [1:0] bus__T_43; // @[OneHot.scala 32:28]
  wire  bus__T_44; // @[CircuitMath.scala 30:8]
  wire [1:0] bus__T_45; // @[Cat.scala 29:58]
  wire  bus__T_48; // @[OneHot.scala 30:18]
  wire [1:0] bus__T_49; // @[OneHot.scala 31:18]
  wire [1:0] bus__GEN_23; // @[OneHot.scala 32:28]
  wire [1:0] bus__T_51; // @[OneHot.scala 32:28]
  wire  bus__T_52; // @[CircuitMath.scala 30:8]
  wire [1:0] bus__T_53; // @[Cat.scala 29:58]
  wire  bus__T_132; // @[Mux.scala 27:72]
  wire  bus__T_133; // @[Mux.scala 27:72]
  wire  bus__T_135; // @[Mux.scala 27:72]
  wire  bus__T_134; // @[Mux.scala 27:72]
  wire  bus_in_0_ar_ready; // @[Mux.scala 27:72]
  reg [2:0] bus__T_59; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_823;
  wire  bus__T_78; // @[Xbar.scala 112:22]
  reg [1:0] bus__T_60; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_824;
  wire  bus__T_77; // @[Xbar.scala 111:75]
  wire  bus__T_79; // @[Xbar.scala 112:34]
  wire  bus__T_80; // @[Xbar.scala 112:80]
  wire  bus__T_82; // @[Xbar.scala 112:48]
  wire  bus_io_in_0_ar_ready; // @[Xbar.scala 130:45]
  wire  bus__T_54; // @[Decoupled.scala 40:37]
  reg  bus__T_302; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_825;
  wire  bus__T_159; // @[Xbar.scala 222:40]
  wire  bus__T_161; // @[Xbar.scala 222:40]
  wire  bus__T_303; // @[Xbar.scala 246:36]
  wire  bus__T_163; // @[Xbar.scala 222:40]
  wire  bus__T_304; // @[Xbar.scala 246:36]
  reg  bus__T_373_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_826;
  wire  bus__T_380; // @[Mux.scala 27:72]
  reg  bus__T_373_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_827;
  wire  bus__T_381; // @[Mux.scala 27:72]
  wire  bus__T_383; // @[Mux.scala 27:72]
  reg  bus__T_373_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_828;
  wire  bus__T_382; // @[Mux.scala 27:72]
  wire  bus__T_384; // @[Mux.scala 27:72]
  wire  bus_in_0_r_valid; // @[Xbar.scala 278:22]
  wire  bus__T_56; // @[Decoupled.scala 40:37]
  wire [2:0] bus__T_306; // @[Cat.scala 29:58]
  reg [2:0] bus__T_313; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_829;
  wire [2:0] bus__T_314; // @[Arbiter.scala 21:30]
  wire [2:0] bus__T_315; // @[Arbiter.scala 21:28]
  wire [5:0] bus__T_316; // @[Cat.scala 29:58]
  wire [4:0] bus__T_317; // @[package.scala 208:48]
  wire [5:0] bus__GEN_24; // @[package.scala 208:43]
  wire [5:0] bus__T_318; // @[package.scala 208:43]
  wire [3:0] bus__T_319; // @[package.scala 208:48]
  wire [5:0] bus__GEN_25; // @[package.scala 208:43]
  wire [5:0] bus__T_320; // @[package.scala 208:43]
  wire [4:0] bus__T_322; // @[Arbiter.scala 22:52]
  wire [5:0] bus__T_323; // @[Arbiter.scala 22:66]
  wire [5:0] bus__GEN_26; // @[Arbiter.scala 22:58]
  wire [5:0] bus__T_324; // @[Arbiter.scala 22:58]
  wire [2:0] bus__T_325; // @[Arbiter.scala 23:29]
  wire [2:0] bus__T_326; // @[Arbiter.scala 23:48]
  wire [2:0] bus__T_327; // @[Arbiter.scala 23:39]
  wire [2:0] bus__T_328; // @[Arbiter.scala 23:18]
  wire  bus__T_340; // @[Xbar.scala 248:69]
  wire  bus__T_344; // @[Xbar.scala 250:63]
  wire  bus__T_374_0; // @[Xbar.scala 262:23]
  wire [35:0] bus__T_389; // @[Mux.scala 27:72]
  wire [35:0] bus__T_390; // @[Mux.scala 27:72]
  wire  bus__T_341; // @[Xbar.scala 248:69]
  wire  bus__T_345; // @[Xbar.scala 250:63]
  wire  bus__T_374_1; // @[Xbar.scala 262:23]
  wire [35:0] bus__T_393; // @[Mux.scala 27:72]
  wire [35:0] bus__T_394; // @[Mux.scala 27:72]
  wire [35:0] bus__T_399; // @[Mux.scala 27:72]
  wire  bus__T_342; // @[Xbar.scala 248:69]
  wire  bus__T_346; // @[Xbar.scala 250:63]
  wire  bus__T_374_2; // @[Xbar.scala 262:23]
  wire [35:0] bus__T_397; // @[Mux.scala 27:72]
  wire [35:0] bus__T_398; // @[Mux.scala 27:72]
  wire [35:0] bus__T_400; // @[Mux.scala 27:72]
  wire  bus_in_0_r_bits_last; // @[Mux.scala 27:72]
  wire  bus__T_58; // @[Xbar.scala 120:45]
  wire [2:0] bus__GEN_27; // @[Xbar.scala 106:30]
  wire [2:0] bus__T_62; // @[Xbar.scala 106:30]
  wire [2:0] bus__GEN_28; // @[Xbar.scala 106:48]
  wire [2:0] bus__T_64; // @[Xbar.scala 106:48]
  wire  bus__T_65; // @[Xbar.scala 107:23]
  wire  bus__T_66; // @[Xbar.scala 107:43]
  wire  bus__T_67; // @[Xbar.scala 107:34]
  wire  bus__T_69; // @[Xbar.scala 107:22]
  wire  bus__T_70; // @[Xbar.scala 107:22]
  wire  bus__T_71; // @[Xbar.scala 108:23]
  wire  bus__T_73; // @[Xbar.scala 108:34]
  wire  bus__T_75; // @[Xbar.scala 108:22]
  wire  bus__T_76; // @[Xbar.scala 108:22]
  wire  bus__T_142; // @[Mux.scala 27:72]
  wire  bus__T_143; // @[Mux.scala 27:72]
  wire  bus__T_145; // @[Mux.scala 27:72]
  wire  bus__T_144; // @[Mux.scala 27:72]
  wire  bus_in_0_aw_ready; // @[Mux.scala 27:72]
  reg  bus__T_113; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_830;
  wire  bus__T_117; // @[Xbar.scala 139:57]
  wire  bus__T_118; // @[Xbar.scala 139:45]
  reg [2:0] bus__T_87; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_831;
  wire  bus__T_106; // @[Xbar.scala 112:22]
  reg [1:0] bus__T_88; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_832;
  wire  bus__T_105; // @[Xbar.scala 111:75]
  wire  bus__T_107; // @[Xbar.scala 112:34]
  wire  bus__T_108; // @[Xbar.scala 112:80]
  wire  bus__T_110; // @[Xbar.scala 112:48]
  wire  bus_io_in_0_aw_ready; // @[Xbar.scala 139:82]
  wire  bus__T_83; // @[Decoupled.scala 40:37]
  reg  bus__T_407; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_833;
  wire  bus__T_165; // @[Xbar.scala 222:40]
  wire  bus__T_167; // @[Xbar.scala 222:40]
  wire  bus__T_408; // @[Xbar.scala 246:36]
  wire  bus__T_169; // @[Xbar.scala 222:40]
  wire  bus__T_409; // @[Xbar.scala 246:36]
  reg  bus__T_478_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_834;
  wire  bus__T_485; // @[Mux.scala 27:72]
  reg  bus__T_478_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_835;
  wire  bus__T_486; // @[Mux.scala 27:72]
  wire  bus__T_488; // @[Mux.scala 27:72]
  reg  bus__T_478_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_836;
  wire  bus__T_487; // @[Mux.scala 27:72]
  wire  bus__T_489; // @[Mux.scala 27:72]
  wire  bus_in_0_b_valid; // @[Xbar.scala 278:22]
  wire  bus__T_85; // @[Decoupled.scala 40:37]
  wire [2:0] bus__GEN_29; // @[Xbar.scala 106:30]
  wire [2:0] bus__T_90; // @[Xbar.scala 106:30]
  wire [2:0] bus__GEN_30; // @[Xbar.scala 106:48]
  wire [2:0] bus__T_92; // @[Xbar.scala 106:48]
  wire  bus__T_93; // @[Xbar.scala 107:23]
  wire  bus__T_94; // @[Xbar.scala 107:43]
  wire  bus__T_95; // @[Xbar.scala 107:34]
  wire  bus__T_97; // @[Xbar.scala 107:22]
  wire  bus__T_98; // @[Xbar.scala 107:22]
  wire  bus__T_99; // @[Xbar.scala 108:23]
  wire  bus__T_101; // @[Xbar.scala 108:34]
  wire  bus__T_103; // @[Xbar.scala 108:22]
  wire  bus__T_104; // @[Xbar.scala 108:22]
  wire  bus_in_0_ar_valid; // @[Xbar.scala 129:45]
  wire  bus__T_115; // @[Xbar.scala 138:45]
  wire  bus_in_0_aw_valid; // @[Xbar.scala 138:82]
  wire  bus__T_120; // @[Xbar.scala 140:54]
  wire  bus__T_122; // @[Decoupled.scala 40:37]
  wire  bus__GEN_2; // @[Xbar.scala 141:38]
  wire  bus__T_123; // @[Decoupled.scala 40:37]
  wire  bus_in_0_w_valid; // @[Xbar.scala 145:43]
  wire  bus__T_152; // @[Mux.scala 27:72]
  wire  bus__T_153; // @[Mux.scala 27:72]
  wire  bus__T_155; // @[Mux.scala 27:72]
  wire  bus__T_154; // @[Mux.scala 27:72]
  wire  bus_in_0_w_ready; // @[Mux.scala 27:72]
  wire  bus__T_126; // @[Xbar.scala 147:50]
  wire  bus_out_0_ar_valid; // @[Xbar.scala 222:40]
  wire  bus_out_1_ar_valid; // @[Xbar.scala 222:40]
  wire  bus_out_2_ar_valid; // @[Xbar.scala 222:40]
  wire  bus_out_0_aw_valid; // @[Xbar.scala 222:40]
  wire  bus_out_1_aw_valid; // @[Xbar.scala 222:40]
  wire  bus_out_2_aw_valid; // @[Xbar.scala 222:40]
  wire  bus__T_176; // @[Xbar.scala 256:60]
  wire  bus__T_182; // @[Xbar.scala 258:23]
  wire  bus__T_184; // @[Xbar.scala 258:12]
  wire  bus__T_185; // @[Xbar.scala 258:12]
  wire  bus__T_197; // @[Xbar.scala 256:60]
  wire  bus__T_203; // @[Xbar.scala 258:23]
  wire  bus__T_205; // @[Xbar.scala 258:12]
  wire  bus__T_206; // @[Xbar.scala 258:12]
  wire  bus__T_220; // @[Xbar.scala 256:60]
  wire  bus__T_226; // @[Xbar.scala 258:23]
  wire  bus__T_228; // @[Xbar.scala 258:12]
  wire  bus__T_229; // @[Xbar.scala 258:12]
  wire  bus__T_241; // @[Xbar.scala 256:60]
  wire  bus__T_247; // @[Xbar.scala 258:23]
  wire  bus__T_249; // @[Xbar.scala 258:12]
  wire  bus__T_250; // @[Xbar.scala 258:12]
  wire  bus__T_264; // @[Xbar.scala 256:60]
  wire  bus__T_270; // @[Xbar.scala 258:23]
  wire  bus__T_272; // @[Xbar.scala 258:12]
  wire  bus__T_273; // @[Xbar.scala 258:12]
  wire  bus__T_285; // @[Xbar.scala 256:60]
  wire  bus__T_291; // @[Xbar.scala 258:23]
  wire  bus__T_293; // @[Xbar.scala 258:12]
  wire  bus__T_294; // @[Xbar.scala 258:12]
  wire  bus__T_329; // @[Arbiter.scala 24:27]
  wire  bus__T_330; // @[Arbiter.scala 24:18]
  wire [2:0] bus__T_331; // @[Arbiter.scala 25:29]
  wire [3:0] bus__T_332; // @[package.scala 199:48]
  wire [2:0] bus__T_333; // @[package.scala 199:53]
  wire [2:0] bus__T_334; // @[package.scala 199:43]
  wire [4:0] bus__T_335; // @[package.scala 199:48]
  wire [2:0] bus__T_336; // @[package.scala 199:53]
  wire [2:0] bus__T_337; // @[package.scala 199:43]
  wire  bus__T_349; // @[Xbar.scala 255:50]
  wire  bus__T_350; // @[Xbar.scala 255:50]
  wire  bus__T_352; // @[Xbar.scala 256:60]
  wire  bus__T_355; // @[Xbar.scala 256:60]
  wire  bus__T_356; // @[Xbar.scala 256:57]
  wire  bus__T_357; // @[Xbar.scala 256:54]
  wire  bus__T_358; // @[Xbar.scala 256:60]
  wire  bus__T_359; // @[Xbar.scala 256:57]
  wire  bus__T_361; // @[Xbar.scala 256:75]
  wire  bus__T_363; // @[Xbar.scala 256:11]
  wire  bus__T_364; // @[Xbar.scala 256:11]
  wire  bus__T_365; // @[Xbar.scala 258:13]
  wire  bus__T_368; // @[Xbar.scala 258:23]
  wire  bus__T_370; // @[Xbar.scala 258:12]
  wire  bus__T_371; // @[Xbar.scala 258:12]
  wire  bus__GEN_17; // @[Xbar.scala 266:21]
  wire  bus__GEN_18; // @[Xbar.scala 267:24]
  wire  bus__T_376_0; // @[Xbar.scala 270:24]
  wire  bus__T_376_1; // @[Xbar.scala 270:24]
  wire  bus__T_376_2; // @[Xbar.scala 270:24]
  wire [2:0] bus__T_411; // @[Cat.scala 29:58]
  reg [2:0] bus__T_418; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_837;
  wire [2:0] bus__T_419; // @[Arbiter.scala 21:30]
  wire [2:0] bus__T_420; // @[Arbiter.scala 21:28]
  wire [5:0] bus__T_421; // @[Cat.scala 29:58]
  wire [4:0] bus__T_422; // @[package.scala 208:48]
  wire [5:0] bus__GEN_31; // @[package.scala 208:43]
  wire [5:0] bus__T_423; // @[package.scala 208:43]
  wire [3:0] bus__T_424; // @[package.scala 208:48]
  wire [5:0] bus__GEN_32; // @[package.scala 208:43]
  wire [5:0] bus__T_425; // @[package.scala 208:43]
  wire [4:0] bus__T_427; // @[Arbiter.scala 22:52]
  wire [5:0] bus__T_428; // @[Arbiter.scala 22:66]
  wire [5:0] bus__GEN_33; // @[Arbiter.scala 22:58]
  wire [5:0] bus__T_429; // @[Arbiter.scala 22:58]
  wire [2:0] bus__T_430; // @[Arbiter.scala 23:29]
  wire [2:0] bus__T_431; // @[Arbiter.scala 23:48]
  wire [2:0] bus__T_432; // @[Arbiter.scala 23:39]
  wire [2:0] bus__T_433; // @[Arbiter.scala 23:18]
  wire  bus__T_434; // @[Arbiter.scala 24:27]
  wire  bus__T_435; // @[Arbiter.scala 24:18]
  wire [2:0] bus__T_436; // @[Arbiter.scala 25:29]
  wire [3:0] bus__T_437; // @[package.scala 199:48]
  wire [2:0] bus__T_438; // @[package.scala 199:53]
  wire [2:0] bus__T_439; // @[package.scala 199:43]
  wire [4:0] bus__T_440; // @[package.scala 199:48]
  wire [2:0] bus__T_441; // @[package.scala 199:53]
  wire [2:0] bus__T_442; // @[package.scala 199:43]
  wire  bus__T_445; // @[Xbar.scala 248:69]
  wire  bus__T_446; // @[Xbar.scala 248:69]
  wire  bus__T_447; // @[Xbar.scala 248:69]
  wire  bus__T_449; // @[Xbar.scala 250:63]
  wire  bus__T_450; // @[Xbar.scala 250:63]
  wire  bus__T_451; // @[Xbar.scala 250:63]
  wire  bus__T_454; // @[Xbar.scala 255:50]
  wire  bus__T_455; // @[Xbar.scala 255:50]
  wire  bus__T_457; // @[Xbar.scala 256:60]
  wire  bus__T_460; // @[Xbar.scala 256:60]
  wire  bus__T_461; // @[Xbar.scala 256:57]
  wire  bus__T_462; // @[Xbar.scala 256:54]
  wire  bus__T_463; // @[Xbar.scala 256:60]
  wire  bus__T_464; // @[Xbar.scala 256:57]
  wire  bus__T_466; // @[Xbar.scala 256:75]
  wire  bus__T_468; // @[Xbar.scala 256:11]
  wire  bus__T_469; // @[Xbar.scala 256:11]
  wire  bus__T_470; // @[Xbar.scala 258:13]
  wire  bus__T_473; // @[Xbar.scala 258:23]
  wire  bus__T_475; // @[Xbar.scala 258:12]
  wire  bus__T_476; // @[Xbar.scala 258:12]
  wire  bus__T_479_0; // @[Xbar.scala 262:23]
  wire  bus__T_479_1; // @[Xbar.scala 262:23]
  wire  bus__T_479_2; // @[Xbar.scala 262:23]
  wire  bus__GEN_20; // @[Xbar.scala 266:21]
  wire  bus__GEN_21; // @[Xbar.scala 267:24]
  wire  bus__T_481_0; // @[Xbar.scala 270:24]
  wire  bus__T_481_1; // @[Xbar.scala 270:24]
  wire  bus__T_481_2; // @[Xbar.scala 270:24]
  wire [2:0] bus__T_492; // @[Mux.scala 27:72]
  wire [2:0] bus__T_493; // @[Mux.scala 27:72]
  wire [2:0] bus__T_494; // @[Mux.scala 27:72]
  wire [2:0] bus__T_495; // @[Mux.scala 27:72]
  wire [2:0] bus__T_496; // @[Mux.scala 27:72]
  wire [2:0] bus__T_497; // @[Mux.scala 27:72]
  wire [2:0] bus__T_498; // @[Mux.scala 27:72]
  wire [2:0] bus__T_499; // @[Mux.scala 27:72]
  wire  converter_auto_in_aw_ready;
  wire  converter_auto_in_aw_valid;
  wire  converter_auto_in_aw_bits_id;
  wire [31:0] converter_auto_in_aw_bits_addr;
  wire  converter_auto_in_w_ready;
  wire  converter_auto_in_w_valid;
  wire [31:0] converter_auto_in_w_bits_data;
  wire [3:0] converter_auto_in_w_bits_strb;
  wire  converter_auto_in_w_bits_last;
  wire  converter_auto_in_b_ready;
  wire  converter_auto_in_b_valid;
  wire [1:0] converter_auto_in_b_bits_resp;
  wire  converter_auto_in_ar_ready;
  wire  converter_auto_in_ar_valid;
  wire  converter_auto_in_ar_bits_id;
  wire [31:0] converter_auto_in_ar_bits_addr;
  wire [2:0] converter_auto_in_ar_bits_size;
  wire  converter_auto_in_r_ready;
  wire  converter_auto_in_r_valid;
  wire [31:0] converter_auto_in_r_bits_data;
  wire [1:0] converter_auto_in_r_bits_resp;
  wire  converter_auto_in_r_bits_last;
  wire  converter_auto_out_aw_ready;
  wire  converter_auto_out_aw_valid;
  wire  converter_auto_out_aw_bits_id;
  wire [29:0] converter_auto_out_aw_bits_addr;
  wire  converter_auto_out_w_ready;
  wire  converter_auto_out_w_valid;
  wire [31:0] converter_auto_out_w_bits_data;
  wire [3:0] converter_auto_out_w_bits_strb;
  wire  converter_auto_out_w_bits_last;
  wire  converter_auto_out_b_ready;
  wire  converter_auto_out_b_valid;
  wire [1:0] converter_auto_out_b_bits_resp;
  wire  converter_auto_out_ar_ready;
  wire  converter_auto_out_ar_valid;
  wire  converter_auto_out_ar_bits_id;
  wire [29:0] converter_auto_out_ar_bits_addr;
  wire [2:0] converter_auto_out_ar_bits_size;
  wire  converter_auto_out_r_ready;
  wire  converter_auto_out_r_valid;
  wire [31:0] converter_auto_out_r_bits_data;
  wire [1:0] converter_auto_out_r_bits_resp;
  wire  converter_auto_out_r_bits_last;
  wire  converter_1_auto_in_ready;
  wire  converter_1_auto_in_valid;
  wire [15:0] converter_1_auto_in_bits_data;
  wire  converter_1_auto_in_bits_last;
  wire  converter_1_auto_out_ready;
  wire  converter_1_auto_out_valid;
  wire [15:0] converter_1_auto_out_bits_data;
  wire  converter_1_auto_out_bits_last;
  wire  converter_2_auto_in_ready;
  wire  converter_2_auto_in_valid;
  wire [7:0] converter_2_auto_in_bits_data;
  wire  converter_2_auto_in_bits_last;
  wire  converter_2_auto_out_ready;
  wire  converter_2_auto_out_valid;
  wire [7:0] converter_2_auto_out_bits_data;
  wire  converter_2_auto_out_bits_last;
  
  assign sram_R0_addr = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_addr;
  assign sram_R0_en   = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_en;
  assign sram_R0_clk  = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_clk;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_data = sram_R0_data;
  assign sram_W0_addr = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_addr;
  assign sram_W0_en   = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_en;
  assign sram_W0_clk  = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_clk;
  assign sram_W0_data = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_data;

  assign widthAdapter__T_4 = widthAdapter_auto_in_valid & widthAdapter_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  assign widthAdapter__T_5 = widthAdapter__T_3 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign widthAdapter__T_6 = widthAdapter__T_3 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign widthAdapter__T_7 = widthAdapter__T_5 ? 3'h0 : widthAdapter__T_6; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign widthAdapter__GEN_0 = widthAdapter__T_4 ? widthAdapter__T_7 : {{1'd0}, widthAdapter__T_3}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign widthAdapter__T_9 = widthAdapter__T_3 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign widthAdapter__T_10 = widthAdapter__T_4 & widthAdapter__T_9; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign widthAdapter__T_12 = widthAdapter__T_3 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign widthAdapter__T_13 = widthAdapter__T_4 & widthAdapter__T_12; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign widthAdapter__T_15 = widthAdapter__T_3 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign widthAdapter__T_16 = widthAdapter__T_4 & widthAdapter__T_15; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign widthAdapter__T_18 = {widthAdapter_auto_in_bits_data,widthAdapter__T_2,widthAdapter__T_1}; // @[Cat.scala 29:58]
  assign widthAdapter_ov0 = widthAdapter__T_5 & widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign widthAdapter__T_25 = widthAdapter__T_23 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign widthAdapter__T_26 = widthAdapter__T_23 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign widthAdapter__T_27 = widthAdapter__T_25 ? 3'h0 : widthAdapter__T_26; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign widthAdapter__GEN_4 = widthAdapter__T_4 ? widthAdapter__T_27 : {{1'd0}, widthAdapter__T_23}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign widthAdapter__T_29 = widthAdapter__T_23 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign widthAdapter__T_30 = widthAdapter__T_4 & widthAdapter__T_29; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign widthAdapter__T_32 = widthAdapter__T_23 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign widthAdapter__T_33 = widthAdapter__T_4 & widthAdapter__T_32; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign widthAdapter__T_35 = widthAdapter__T_23 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign widthAdapter__T_36 = widthAdapter__T_4 & widthAdapter__T_35; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign widthAdapter__T_39 = {widthAdapter_auto_in_bits_last,widthAdapter__T_22,widthAdapter__T_21,widthAdapter__T_20}; // @[Cat.scala 29:58]
  assign widthAdapter_ov1 = widthAdapter__T_25 & widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign widthAdapter__T_46 = widthAdapter__T_44 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign widthAdapter__T_47 = widthAdapter__T_44 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign widthAdapter__T_48 = widthAdapter__T_46 ? 3'h0 : widthAdapter__T_47; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign widthAdapter__GEN_8 = widthAdapter__T_4 ? widthAdapter__T_48 : {{1'd0}, widthAdapter__T_44}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign widthAdapter_ov2 = widthAdapter__T_46 & widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign widthAdapter__T_66 = widthAdapter__T_64 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign widthAdapter__T_67 = widthAdapter__T_64 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign widthAdapter__T_68 = widthAdapter__T_66 ? 3'h0 : widthAdapter__T_67; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign widthAdapter__GEN_12 = widthAdapter__T_4 ? widthAdapter__T_68 : {{1'd0}, widthAdapter__T_64}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign widthAdapter_ov3 = widthAdapter__T_66 & widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign widthAdapter__T_86 = widthAdapter__T_84 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign widthAdapter__T_87 = widthAdapter__T_84 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign widthAdapter__T_88 = widthAdapter__T_86 ? 3'h0 : widthAdapter__T_87; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign widthAdapter__GEN_16 = widthAdapter__T_4 ? widthAdapter__T_88 : {{1'd0}, widthAdapter__T_84}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign widthAdapter_ov4 = widthAdapter__T_86 & widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign widthAdapter__T_101 = widthAdapter_ov0 == widthAdapter_ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  assign widthAdapter__T_103 = widthAdapter__T_101 | widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign widthAdapter__T_104 = ~widthAdapter__T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign widthAdapter__T_105 = widthAdapter_ov0 == widthAdapter_ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  assign widthAdapter__T_107 = widthAdapter__T_105 | widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign widthAdapter__T_108 = ~widthAdapter__T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign widthAdapter__T_109 = widthAdapter_ov0 == widthAdapter_ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  assign widthAdapter__T_111 = widthAdapter__T_109 | widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign widthAdapter__T_112 = ~widthAdapter__T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign widthAdapter__T_113 = widthAdapter_ov0 == widthAdapter_ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  assign widthAdapter__T_115 = widthAdapter__T_113 | widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign widthAdapter__T_116 = ~widthAdapter__T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign widthAdapter_auto_in_ready = widthAdapter_auto_out_ready; // @[LazyModule.scala 173:31]
  assign widthAdapter_auto_out_valid = widthAdapter__T_5 & widthAdapter_auto_in_valid; // @[LazyModule.scala 173:49]
  assign widthAdapter_auto_out_bits_data = {widthAdapter__T_18,widthAdapter__T}; // @[LazyModule.scala 173:49]
  assign widthAdapter_auto_out_bits_last = widthAdapter__T_39 != 4'h0; // @[LazyModule.scala 173:49]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_load_input = fft_fft_SDFChainRadix22_sdf_stages_0_io_cntr < 9'h1; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_0_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_0_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_47 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_49 = fft_fft_SDFChainRadix22_sdf_stages_0__T_47[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_52 = $signed(fft_fft_SDFChainRadix22_sdf_stages_0__T_49) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_0__T_52[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_0_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_0_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_54 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_56 = fft_fft_SDFChainRadix22_sdf_stages_0__T_54[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_59 = $signed(fft_fft_SDFChainRadix22_sdf_stages_0__T_56) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_0__T_59[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_0_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_0_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_0_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_0_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_30 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_32 = fft_fft_SDFChainRadix22_sdf_stages_0__T_30[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_35 = $signed(fft_fft_SDFChainRadix22_sdf_stages_0__T_32) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_0__T_35[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_37 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_0_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_39 = fft_fft_SDFChainRadix22_sdf_stages_0__T_37[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_0__T_42 = $signed(fft_fft_SDFChainRadix22_sdf_stages_0__T_39) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_0__T_42[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_0_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_0_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_0_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_0_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_0_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_0_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_load_input = fft_fft_SDFChainRadix22_sdf_stages_1_io_cntr < 9'h2; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_1_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_1_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_50 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_52 = fft_fft_SDFChainRadix22_sdf_stages_1__T_50[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_55 = $signed(fft_fft_SDFChainRadix22_sdf_stages_1__T_52) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_1__T_55[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_1_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_1_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_57 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_59 = fft_fft_SDFChainRadix22_sdf_stages_1__T_57[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_62 = $signed(fft_fft_SDFChainRadix22_sdf_stages_1__T_59) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_1__T_62[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_1_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_1_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_1_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_1_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_33 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_35 = fft_fft_SDFChainRadix22_sdf_stages_1__T_33[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_38 = $signed(fft_fft_SDFChainRadix22_sdf_stages_1__T_35) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_1__T_38[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_40 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_1_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_42 = fft_fft_SDFChainRadix22_sdf_stages_1__T_40[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_1__T_45 = $signed(fft_fft_SDFChainRadix22_sdf_stages_1__T_42) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_1__T_45[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_1_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_1_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_1_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_1_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_1_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_1_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_load_input = fft_fft_SDFChainRadix22_sdf_stages_2_io_cntr < 9'h4; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_2_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_2_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_56 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_58 = fft_fft_SDFChainRadix22_sdf_stages_2__T_56[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_61 = $signed(fft_fft_SDFChainRadix22_sdf_stages_2__T_58) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_2__T_61[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_2_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_2_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_63 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_65 = fft_fft_SDFChainRadix22_sdf_stages_2__T_63[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_68 = $signed(fft_fft_SDFChainRadix22_sdf_stages_2__T_65) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_2__T_68[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_2_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_2_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_2_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_2_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_39 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_41 = fft_fft_SDFChainRadix22_sdf_stages_2__T_39[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_44 = $signed(fft_fft_SDFChainRadix22_sdf_stages_2__T_41) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_2__T_44[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_46 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_2_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_48 = fft_fft_SDFChainRadix22_sdf_stages_2__T_46[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_2__T_51 = $signed(fft_fft_SDFChainRadix22_sdf_stages_2__T_48) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_2__T_51[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_2_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_2_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_2_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_2_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_2_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_2_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_load_input = fft_fft_SDFChainRadix22_sdf_stages_3_io_cntr < 9'h8; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_3_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_3_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_68 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_70 = fft_fft_SDFChainRadix22_sdf_stages_3__T_68[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_73 = $signed(fft_fft_SDFChainRadix22_sdf_stages_3__T_70) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_3__T_73[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_3_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_3_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_75 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_77 = fft_fft_SDFChainRadix22_sdf_stages_3__T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_80 = $signed(fft_fft_SDFChainRadix22_sdf_stages_3__T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_3__T_80[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_3_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_3_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_3_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_3_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_51 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_53 = fft_fft_SDFChainRadix22_sdf_stages_3__T_51[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_56 = $signed(fft_fft_SDFChainRadix22_sdf_stages_3__T_53) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_3__T_56[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_58 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_3_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_60 = fft_fft_SDFChainRadix22_sdf_stages_3__T_58[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_3__T_63 = $signed(fft_fft_SDFChainRadix22_sdf_stages_3__T_60) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_3__T_63[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_3_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_3_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_3_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_3_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_3_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_3_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_load_input = fft_fft_SDFChainRadix22_sdf_stages_4_io_cntr < 9'h10; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_4_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_4_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_92 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_94 = fft_fft_SDFChainRadix22_sdf_stages_4__T_92[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_97 = $signed(fft_fft_SDFChainRadix22_sdf_stages_4__T_94) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_4__T_97[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_4_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_4_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_99 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_101 = fft_fft_SDFChainRadix22_sdf_stages_4__T_99[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_104 = $signed(fft_fft_SDFChainRadix22_sdf_stages_4__T_101) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_4__T_104[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_4_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_4_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_4_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_4_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_75 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_77 = fft_fft_SDFChainRadix22_sdf_stages_4__T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_80 = $signed(fft_fft_SDFChainRadix22_sdf_stages_4__T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_4__T_80[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_82 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_4_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_84 = fft_fft_SDFChainRadix22_sdf_stages_4__T_82[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_4__T_87 = $signed(fft_fft_SDFChainRadix22_sdf_stages_4__T_84) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_4__T_87[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_4_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_4_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_4_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_4_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_4_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_4_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_load_input = fft_fft_SDFChainRadix22_sdf_stages_5_io_cntr < 9'h20; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_5_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_5_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_140 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_142 = fft_fft_SDFChainRadix22_sdf_stages_5__T_140[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_145 = $signed(fft_fft_SDFChainRadix22_sdf_stages_5__T_142) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_5__T_145[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_5_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_5_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_147 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_149 = fft_fft_SDFChainRadix22_sdf_stages_5__T_147[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_152 = $signed(fft_fft_SDFChainRadix22_sdf_stages_5__T_149) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_5__T_152[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_5_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_5_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_5_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_5_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_123 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_125 = fft_fft_SDFChainRadix22_sdf_stages_5__T_123[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_128 = $signed(fft_fft_SDFChainRadix22_sdf_stages_5__T_125) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_5__T_128[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_130 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_5_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_132 = fft_fft_SDFChainRadix22_sdf_stages_5__T_130[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_5__T_135 = $signed(fft_fft_SDFChainRadix22_sdf_stages_5__T_132) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_5__T_135[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_5_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_5_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_5_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_5_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_5_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_5_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_load_input = fft_fft_SDFChainRadix22_sdf_stages_6_io_cntr < 9'h40; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_6_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_6_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_236 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_238 = fft_fft_SDFChainRadix22_sdf_stages_6__T_236[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_241 = $signed(fft_fft_SDFChainRadix22_sdf_stages_6__T_238) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_6__T_241[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_6_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_6_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_243 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_245 = fft_fft_SDFChainRadix22_sdf_stages_6__T_243[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_248 = $signed(fft_fft_SDFChainRadix22_sdf_stages_6__T_245) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_6__T_248[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_6_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_6_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_6_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_6_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_219 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_221 = fft_fft_SDFChainRadix22_sdf_stages_6__T_219[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_224 = $signed(fft_fft_SDFChainRadix22_sdf_stages_6__T_221) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_6__T_224[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_226 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_6_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_228 = fft_fft_SDFChainRadix22_sdf_stages_6__T_226[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_6__T_231 = $signed(fft_fft_SDFChainRadix22_sdf_stages_6__T_228) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_6__T_231[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_6_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_6_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_6_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_6_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_6_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_6_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_load_input = fft_fft_SDFChainRadix22_sdf_stages_7_io_cntr < 9'h80; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_7_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_7_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_428 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_430 = fft_fft_SDFChainRadix22_sdf_stages_7__T_428[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_433 = $signed(fft_fft_SDFChainRadix22_sdf_stages_7__T_430) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_7__T_433[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_7_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_7_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_435 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_437 = fft_fft_SDFChainRadix22_sdf_stages_7__T_435[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_440 = $signed(fft_fft_SDFChainRadix22_sdf_stages_7__T_437) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_7__T_440[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_7_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_7_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_7_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_7_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_411 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_413 = fft_fft_SDFChainRadix22_sdf_stages_7__T_411[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_416 = $signed(fft_fft_SDFChainRadix22_sdf_stages_7__T_413) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_7__T_416[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_418 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_7_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_420 = fft_fft_SDFChainRadix22_sdf_stages_7__T_418[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_7__T_423 = $signed(fft_fft_SDFChainRadix22_sdf_stages_7__T_420) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_7__T_423[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_7_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_7_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_7_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_7_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_7_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_7_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_clk = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_clk;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_en = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_en;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_addr = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_addr;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_data_imag = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_data[15:0];
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_data_real = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_R0_data[31:16];
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_clk = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_clk;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_en = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_en;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_addr = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_addr;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_SRAM_depth_256_width_32_mem_ext_W0_data = {fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_data_real,fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_data_imag};
  assign fft_fft_SDFChainRadix22_sdf_stages_8_load_input = fft_fft_SDFChainRadix22_sdf_stages_8_io_cntr < 9'h100; // @[UIntTypeClass.scala 52:47]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_feedback_real = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_data_real; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_1_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_8_feedback_real) - $signed(fft_fft_SDFChainRadix22_sdf_stages_8_io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_57 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_59 = fft_fft_SDFChainRadix22_sdf_stages_8__T_57[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_62 = $signed(fft_fft_SDFChainRadix22_sdf_stages_8__T_59) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butterfly_outputs_1_real = fft_fft_SDFChainRadix22_sdf_stages_8__T_62[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_feedback_imag = fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_data_imag; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_1_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_8_feedback_imag) - $signed(fft_fft_SDFChainRadix22_sdf_stages_8_io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_64 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_66 = fft_fft_SDFChainRadix22_sdf_stages_8__T_64[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_69 = $signed(fft_fft_SDFChainRadix22_sdf_stages_8__T_66) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butterfly_outputs_1_imag = fft_fft_SDFChainRadix22_sdf_stages_8__T_69[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_22 = fft_fft_SDFChainRadix22_sdf_stages_8_value + 8'h1; // @[Counter.scala 39:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_0_real = $signed(fft_fft_SDFChainRadix22_sdf_stages_8_feedback_real) + $signed(fft_fft_SDFChainRadix22_sdf_stages_8_io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_0_imag = $signed(fft_fft_SDFChainRadix22_sdf_stages_8_feedback_imag) + $signed(fft_fft_SDFChainRadix22_sdf_stages_8_io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_40 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_42 = fft_fft_SDFChainRadix22_sdf_stages_8__T_40[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_45 = $signed(fft_fft_SDFChainRadix22_sdf_stages_8__T_42) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butt_out_0_real = fft_fft_SDFChainRadix22_sdf_stages_8__T_45[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_47 = {$signed(fft_fft_SDFChainRadix22_sdf_stages_8_butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_49 = fft_fft_SDFChainRadix22_sdf_stages_8__T_47[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_8__T_52 = $signed(fft_fft_SDFChainRadix22_sdf_stages_8__T_49) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_butt_out_0_imag = fft_fft_SDFChainRadix22_sdf_stages_8__T_52[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_io_out_real = fft_fft_SDFChainRadix22_sdf_stages_8_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_8_feedback_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_8_butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_io_out_imag = fft_fft_SDFChainRadix22_sdf_stages_8_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_8_feedback_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_8_butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_addr = fft_fft_SDFChainRadix22_sdf_stages_8_value; // @[ShiftRegisterMem.scala 53:25]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_en = fft_fft_SDFChainRadix22_sdf_stages_8_io_en; // @[ShiftRegisterMem.scala 48:28 Counter.scala 39:13]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_R0_clk = fft_fft_SDFChainRadix22_sdf_stages_8_clock; // @[ShiftRegisterMem.scala 53:25]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_addr = fft_fft_SDFChainRadix22_sdf_stages_8__T_26;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_en = fft_fft_SDFChainRadix22_sdf_stages_8_io_en; // @[ShiftRegisterMem.scala 48:28]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_clk = fft_fft_SDFChainRadix22_sdf_stages_8_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_data_real = fft_fft_SDFChainRadix22_sdf_stages_8_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_8_io_in_real) : $signed(fft_fft_SDFChainRadix22_sdf_stages_8_butterfly_outputs_1_real);
  assign fft_fft_SDFChainRadix22_sdf_stages_8_SRAM_depth_256_width_32_mem_W0_data_imag = fft_fft_SDFChainRadix22_sdf_stages_8_load_input ? $signed(fft_fft_SDFChainRadix22_sdf_stages_8_io_in_imag) : $signed(fft_fft_SDFChainRadix22_sdf_stages_8_butterfly_outputs_1_imag);
  assign fft_fft_SDFChainRadix22__T_46 = fft_fft_SDFChainRadix22_io_in_ready & fft_fft_SDFChainRadix22_io_in_valid; // @[Decoupled.scala 40:37]
  assign fft_fft_SDFChainRadix22_fireLast = fft_fft_SDFChainRadix22_io_lastIn & fft_fft_SDFChainRadix22__T_46; // @[SDFChainRadix22.scala 79:28]
  assign fft_fft_SDFChainRadix22__T_48 = 9'h9 - 9'h1; // @[SDFChainRadix22.scala 81:45]
  assign fft_fft_SDFChainRadix22__T_49 = fft_fft_SDFChainRadix22__T_48[3:0];
  assign fft_fft_SDFChainRadix22__T_53 = 2'h0 == fft_fft_SDFChainRadix22_state; // @[Conditional.scala 37:30]
  assign fft_fft_SDFChainRadix22__GEN_0 = fft_fft_SDFChainRadix22__T_46 ? 2'h1 : fft_fft_SDFChainRadix22_state; // @[SDFChainRadix22.scala 90:27]
  assign fft_fft_SDFChainRadix22__T_56 = 2'h1 == fft_fft_SDFChainRadix22_state; // @[Conditional.scala 37:30]
  assign fft_fft_SDFChainRadix22__GEN_1 = fft_fft_SDFChainRadix22_fireLast ? 2'h2 : fft_fft_SDFChainRadix22_state; // @[SDFChainRadix22.scala 93:23]
  assign fft_fft_SDFChainRadix22__T_57 = 2'h2 == fft_fft_SDFChainRadix22_state; // @[Conditional.scala 37:30]
  assign fft_fft_SDFChainRadix22__GEN_2 = fft_fft_SDFChainRadix22_io_lastOut ? 2'h0 : fft_fft_SDFChainRadix22_state; // @[SDFChainRadix22.scala 98:25]
  assign fft_fft_SDFChainRadix22__GEN_3 = fft_fft_SDFChainRadix22__T_57 ? fft_fft_SDFChainRadix22__GEN_2 : fft_fft_SDFChainRadix22_state; // @[Conditional.scala 39:67]
  assign fft_fft_SDFChainRadix22__GEN_4 = fft_fft_SDFChainRadix22__T_56 ? fft_fft_SDFChainRadix22__GEN_1 : fft_fft_SDFChainRadix22__GEN_3; // @[Conditional.scala 39:67]
  assign fft_fft_SDFChainRadix22_state_next = fft_fft_SDFChainRadix22__T_53 ? fft_fft_SDFChainRadix22__GEN_0 : fft_fft_SDFChainRadix22__GEN_4; // @[Conditional.scala 40:58]
  assign fft_fft_SDFChainRadix22__T_59 = 10'h200 - 10'h1; // @[SDFChainRadix22.scala 111:44]
  assign fft_fft_SDFChainRadix22__GEN_2109 = {{1'd0}, fft_fft_SDFChainRadix22_cntValidOut}; // @[SDFChainRadix22.scala 111:29]
  assign fft_fft_SDFChainRadix22__T_60 = fft_fft_SDFChainRadix22__GEN_2109 == fft_fft_SDFChainRadix22__T_59; // @[SDFChainRadix22.scala 111:29]
  assign fft_fft_SDFChainRadix22__T_61 = fft_fft_SDFChainRadix22_io_out_ready & fft_fft_SDFChainRadix22_io_out_valid; // @[Decoupled.scala 40:37]
  assign fft_fft_SDFChainRadix22_pktEnd = fft_fft_SDFChainRadix22__T_60 & fft_fft_SDFChainRadix22__T_61; // @[SDFChainRadix22.scala 111:52]
  assign fft_fft_SDFChainRadix22__T_62 = fft_fft_SDFChainRadix22_state_next == 2'h0; // @[SDFChainRadix22.scala 114:20]
  assign fft_fft_SDFChainRadix22_cntr_wires_0 = fft_fft_SDFChainRadix22_cnt[8:0]; // @[SDFChainRadix22.scala 52:24 SDFChainRadix22.scala 185:29]
  assign fft_fft_SDFChainRadix22__GEN_20 = 4'h1 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22_cntr_wires_0; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_21 = 4'h2 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22__GEN_20; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_22 = 4'h3 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22__GEN_21; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_23 = 4'h4 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22__GEN_22; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_24 = 4'h5 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22__GEN_23; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_25 = 4'h6 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22__GEN_24; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_26 = 4'h7 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22__GEN_25; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_27 = 4'h8 == fft_fft_SDFChainRadix22__T_49 ? fft_fft_SDFChainRadix22_cntr_wires_0 : fft_fft_SDFChainRadix22__GEN_26; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__GEN_2110 = {{1'd0}, fft_fft_SDFChainRadix22__GEN_27}; // @[SDFChainRadix22.scala 126:79]
  assign fft_fft_SDFChainRadix22__T_76 = fft_fft_SDFChainRadix22__T_62 & fft_fft_SDFChainRadix22_pktEnd; // @[SDFChainRadix22.scala 130:31]
  assign fft_fft_SDFChainRadix22__T_77 = fft_fft_SDFChainRadix22__T_76 | fft_fft_SDFChainRadix22_pktEnd; // @[SDFChainRadix22.scala 130:42]
  assign fft_fft_SDFChainRadix22__T_80 = fft_fft_SDFChainRadix22_cntValidOut + 9'h1; // @[SDFChainRadix22.scala 134:32]
  assign fft_fft_SDFChainRadix22__T_83 = fft_fft_SDFChainRadix22_state == 2'h2; // @[SDFChainRadix22.scala 144:90]
  assign fft_fft_SDFChainRadix22__T_122 = fft_fft_SDFChainRadix22__T_83 & fft_fft_SDFChainRadix22_io_out_ready; // @[SDFChainRadix22.scala 173:54]
  assign fft_fft_SDFChainRadix22_enableInit = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 173:33]
  assign fft_fft_SDFChainRadix22__T_125 = fft_fft_SDFChainRadix22_cnt + 10'h1; // @[SDFChainRadix22.scala 179:16]
  assign fft_fft_SDFChainRadix22__T_145 = 10'h200 - 10'h2; // @[SDFChainRadix22.scala 193:37]
  assign fft_fft_SDFChainRadix22__T_146 = fft_fft_SDFChainRadix22__GEN_2110 == fft_fft_SDFChainRadix22__T_145; // @[SDFChainRadix22.scala 193:22]
  assign fft_fft_SDFChainRadix22__T_147 = fft_fft_SDFChainRadix22__T_146 & fft_fft_SDFChainRadix22_enableInit; // @[SDFChainRadix22.scala 193:44]
  assign fft_fft_SDFChainRadix22__GEN_45 = fft_fft_SDFChainRadix22__T_62 ? 1'h0 : fft_fft_SDFChainRadix22_initialOutDone; // @[SDFChainRadix22.scala 196:36]
  assign fft_fft_SDFChainRadix22__GEN_46 = fft_fft_SDFChainRadix22__T_147 | fft_fft_SDFChainRadix22__GEN_45; // @[SDFChainRadix22.scala 193:60]
  assign fft_fft_SDFChainRadix22__T_166 = fft_fft_SDFChainRadix22_cntr_wires_0 - 9'h0; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_167 = fft_fft_SDFChainRadix22__T_166[0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_171 = 9'h1 - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_173 = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_171; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_174 = fft_fft_SDFChainRadix22__T_173[1:0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_178 = 9'h3 - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_180 = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_178; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_181 = fft_fft_SDFChainRadix22__T_180[2:0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_185 = 9'h7 - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_187 = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_185; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_188 = fft_fft_SDFChainRadix22__T_187[3:0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_192 = 9'hf - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_194 = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_192; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_195 = fft_fft_SDFChainRadix22__T_194[4:0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_199 = 9'h1f - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_201 = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_199; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_202 = fft_fft_SDFChainRadix22__T_201[5:0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_206 = 9'h3f - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_208 = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_206; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_209 = fft_fft_SDFChainRadix22__T_208[6:0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_213 = 9'h7f - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_215 = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_213; // @[SDFChainRadix22.scala 224:38]
  assign fft_fft_SDFChainRadix22__T_216 = fft_fft_SDFChainRadix22__T_215[7:0]; // @[SDFChainRadix22.scala 224:92]
  assign fft_fft_SDFChainRadix22__T_220 = 9'hff - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign fft_fft_SDFChainRadix22__T_255 = fft_fft_SDFChainRadix22__T_173[2:0];
  assign fft_fft_SDFChainRadix22__GEN_52 = 3'h3 == fft_fft_SDFChainRadix22__T_255 ? 2'h2 : 2'h0; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_53 = 3'h4 == fft_fft_SDFChainRadix22__T_255 ? 2'h0 : fft_fft_SDFChainRadix22__GEN_52; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_54 = 3'h5 == fft_fft_SDFChainRadix22__T_255 ? 2'h1 : fft_fft_SDFChainRadix22__GEN_53; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_55 = 3'h6 == fft_fft_SDFChainRadix22__T_255 ? 2'h0 : fft_fft_SDFChainRadix22__GEN_54; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_56 = 3'h7 == fft_fft_SDFChainRadix22__T_255 ? 2'h3 : fft_fft_SDFChainRadix22__GEN_55; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_59 = 2'h1 == fft_fft_SDFChainRadix22__GEN_56 ? $signed(16'sh2d41) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_60 = 2'h1 == fft_fft_SDFChainRadix22__GEN_56 ? $signed(-16'sh2d41) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_61 = 2'h2 == fft_fft_SDFChainRadix22__GEN_56 ? $signed(16'sh0) : $signed(fft_fft_SDFChainRadix22__GEN_59); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_62 = 2'h2 == fft_fft_SDFChainRadix22__GEN_56 ? $signed(-16'sh4000) : $signed(fft_fft_SDFChainRadix22__GEN_60); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_63 = 2'h3 == fft_fft_SDFChainRadix22__GEN_56 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_61); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22_twiddles_1_imag = 2'h3 == fft_fft_SDFChainRadix22__GEN_56 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_62); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__T_261 = $signed(fft_fft_SDFChainRadix22__GEN_63) + $signed(fft_fft_SDFChainRadix22_twiddles_1_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_outputWires_0_real = fft_fft_SDFChainRadix22_sdf_stages_0_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  assign fft_fft_SDFChainRadix22_outputWires_0_imag = fft_fft_SDFChainRadix22_sdf_stages_0_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  assign fft_fft_SDFChainRadix22__T_262 = $signed(fft_fft_SDFChainRadix22_outputWires_0_real) + $signed(fft_fft_SDFChainRadix22_outputWires_0_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_263 = $signed(fft_fft_SDFChainRadix22_outputWires_0_imag) - $signed(fft_fft_SDFChainRadix22_outputWires_0_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__GEN_2112 = {{1{fft_fft_SDFChainRadix22_outputWires_0_real[15]}},fft_fft_SDFChainRadix22_outputWires_0_real}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_264 = $signed(fft_fft_SDFChainRadix22__GEN_2112) * $signed(fft_fft_SDFChainRadix22__T_261); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2113 = {{1{fft_fft_SDFChainRadix22_twiddles_1_imag[15]}},fft_fft_SDFChainRadix22_twiddles_1_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_265 = $signed(fft_fft_SDFChainRadix22__T_262) * $signed(fft_fft_SDFChainRadix22__GEN_2113); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2114 = {{1{fft_fft_SDFChainRadix22__GEN_63[15]}},fft_fft_SDFChainRadix22__GEN_63}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_266 = $signed(fft_fft_SDFChainRadix22__T_263) * $signed(fft_fft_SDFChainRadix22__GEN_2114); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_267 = $signed(fft_fft_SDFChainRadix22__T_264) - $signed(fft_fft_SDFChainRadix22__T_265); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__T_268 = $signed(fft_fft_SDFChainRadix22__T_264) + $signed(fft_fft_SDFChainRadix22__T_266); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_274 = $signed(fft_fft_SDFChainRadix22__T_267) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_275 = fft_fft_SDFChainRadix22__T_274[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_278 = $signed(fft_fft_SDFChainRadix22__T_268) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_279 = fft_fft_SDFChainRadix22__T_278[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_286 = fft_fft_SDFChainRadix22_sdf_stages_2_io_cntr < 9'h4; // @[SDFChainRadix22.scala 328:32]
  assign fft_fft_SDFChainRadix22__T_287 = fft_fft_SDFChainRadix22_sdf_stages_2_io_cntr < 9'h6; // @[SDFChainRadix22.scala 328:78]
  assign fft_fft_SDFChainRadix22__T_288 = fft_fft_SDFChainRadix22__T_287 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign fft_fft_SDFChainRadix22__T_289 = fft_fft_SDFChainRadix22__T_286 ? 1'h0 : fft_fft_SDFChainRadix22__T_288; // @[SDFChainRadix22.scala 328:19]
  assign fft_fft_SDFChainRadix22_outputWires_1_real = fft_fft_SDFChainRadix22_sdf_stages_1_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__T_295 = 16'sh0 - $signed(fft_fft_SDFChainRadix22_outputWires_1_real); // @[FixedPointTypeClass.scala 39:43]
  assign fft_fft_SDFChainRadix22_outputWires_1_imag = fft_fft_SDFChainRadix22_sdf_stages_1_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__T_387 = fft_fft_SDFChainRadix22__T_187[4:0];
  assign fft_fft_SDFChainRadix22__GEN_82 = 5'h9 == fft_fft_SDFChainRadix22__T_387 ? 4'h2 : 4'h0; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_83 = 5'ha == fft_fft_SDFChainRadix22__T_387 ? 4'h4 : fft_fft_SDFChainRadix22__GEN_82; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_84 = 5'hb == fft_fft_SDFChainRadix22__T_387 ? 4'h6 : fft_fft_SDFChainRadix22__GEN_83; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_85 = 5'hc == fft_fft_SDFChainRadix22__T_387 ? 4'h8 : fft_fft_SDFChainRadix22__GEN_84; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_86 = 5'hd == fft_fft_SDFChainRadix22__T_387 ? 4'ha : fft_fft_SDFChainRadix22__GEN_85; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_87 = 5'he == fft_fft_SDFChainRadix22__T_387 ? 4'hb : fft_fft_SDFChainRadix22__GEN_86; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_88 = 5'hf == fft_fft_SDFChainRadix22__T_387 ? 4'hc : fft_fft_SDFChainRadix22__GEN_87; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_89 = 5'h10 == fft_fft_SDFChainRadix22__T_387 ? 4'h0 : fft_fft_SDFChainRadix22__GEN_88; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_90 = 5'h11 == fft_fft_SDFChainRadix22__T_387 ? 4'h1 : fft_fft_SDFChainRadix22__GEN_89; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_91 = 5'h12 == fft_fft_SDFChainRadix22__T_387 ? 4'h2 : fft_fft_SDFChainRadix22__GEN_90; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_92 = 5'h13 == fft_fft_SDFChainRadix22__T_387 ? 4'h3 : fft_fft_SDFChainRadix22__GEN_91; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_93 = 5'h14 == fft_fft_SDFChainRadix22__T_387 ? 4'h4 : fft_fft_SDFChainRadix22__GEN_92; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_94 = 5'h15 == fft_fft_SDFChainRadix22__T_387 ? 4'h5 : fft_fft_SDFChainRadix22__GEN_93; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_95 = 5'h16 == fft_fft_SDFChainRadix22__T_387 ? 4'h6 : fft_fft_SDFChainRadix22__GEN_94; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_96 = 5'h17 == fft_fft_SDFChainRadix22__T_387 ? 4'h7 : fft_fft_SDFChainRadix22__GEN_95; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_97 = 5'h18 == fft_fft_SDFChainRadix22__T_387 ? 4'h0 : fft_fft_SDFChainRadix22__GEN_96; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_98 = 5'h19 == fft_fft_SDFChainRadix22__T_387 ? 4'h3 : fft_fft_SDFChainRadix22__GEN_97; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_99 = 5'h1a == fft_fft_SDFChainRadix22__T_387 ? 4'h6 : fft_fft_SDFChainRadix22__GEN_98; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_100 = 5'h1b == fft_fft_SDFChainRadix22__T_387 ? 4'h9 : fft_fft_SDFChainRadix22__GEN_99; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_101 = 5'h1c == fft_fft_SDFChainRadix22__T_387 ? 4'hb : fft_fft_SDFChainRadix22__GEN_100; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_102 = 5'h1d == fft_fft_SDFChainRadix22__T_387 ? 4'hd : fft_fft_SDFChainRadix22__GEN_101; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_103 = 5'h1e == fft_fft_SDFChainRadix22__T_387 ? 4'he : fft_fft_SDFChainRadix22__GEN_102; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_104 = 5'h1f == fft_fft_SDFChainRadix22__T_387 ? 4'hf : fft_fft_SDFChainRadix22__GEN_103; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_107 = 4'h1 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh3ec5) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_108 = 4'h1 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'shc7c) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_109 = 4'h2 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_107); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_110 = 4'h2 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_108); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_111 = 4'h3 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_109); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_112 = 4'h3 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_110); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_113 = 4'h4 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_111); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_114 = 4'h4 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_112); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_115 = 4'h5 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_113); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_116 = 4'h5 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_114); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_117 = 4'h6 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_115); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_118 = 4'h6 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_116); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_119 = 4'h7 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_117); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_120 = 4'h7 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_118); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_121 = 4'h8 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh0) : $signed(fft_fft_SDFChainRadix22__GEN_119); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_122 = 4'h8 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh4000) : $signed(fft_fft_SDFChainRadix22__GEN_120); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_123 = 4'h9 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_121); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_124 = 4'h9 == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_122); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_125 = 4'ha == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_123); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_126 = 4'ha == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_124); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_127 = 4'hb == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_125); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_128 = 4'hb == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_126); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_129 = 4'hc == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_127); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_130 = 4'hc == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_128); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_131 = 4'hd == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_129); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_132 = 4'hd == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_130); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_133 = 4'he == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_131); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_134 = 4'he == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_132); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_135 = 4'hf == fft_fft_SDFChainRadix22__GEN_104 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_133); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22_twiddles_3_imag = 4'hf == fft_fft_SDFChainRadix22__GEN_104 ? $signed(16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_134); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__T_393 = $signed(fft_fft_SDFChainRadix22__GEN_135) + $signed(fft_fft_SDFChainRadix22_twiddles_3_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_outputWires_2_real = fft_fft_SDFChainRadix22_sdf_stages_2_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22_outputWires_2_imag = fft_fft_SDFChainRadix22_sdf_stages_2_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22__T_394 = $signed(fft_fft_SDFChainRadix22_outputWires_2_real) + $signed(fft_fft_SDFChainRadix22_outputWires_2_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_395 = $signed(fft_fft_SDFChainRadix22_outputWires_2_imag) - $signed(fft_fft_SDFChainRadix22_outputWires_2_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__GEN_2115 = {{1{fft_fft_SDFChainRadix22_outputWires_2_real[15]}},fft_fft_SDFChainRadix22_outputWires_2_real}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_396 = $signed(fft_fft_SDFChainRadix22__GEN_2115) * $signed(fft_fft_SDFChainRadix22__T_393); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2116 = {{1{fft_fft_SDFChainRadix22_twiddles_3_imag[15]}},fft_fft_SDFChainRadix22_twiddles_3_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_397 = $signed(fft_fft_SDFChainRadix22__T_394) * $signed(fft_fft_SDFChainRadix22__GEN_2116); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2117 = {{1{fft_fft_SDFChainRadix22__GEN_135[15]}},fft_fft_SDFChainRadix22__GEN_135}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_398 = $signed(fft_fft_SDFChainRadix22__T_395) * $signed(fft_fft_SDFChainRadix22__GEN_2117); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_399 = $signed(fft_fft_SDFChainRadix22__T_396) - $signed(fft_fft_SDFChainRadix22__T_397); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__T_400 = $signed(fft_fft_SDFChainRadix22__T_396) + $signed(fft_fft_SDFChainRadix22__T_398); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_406 = $signed(fft_fft_SDFChainRadix22__T_399) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_407 = fft_fft_SDFChainRadix22__T_406[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_410 = $signed(fft_fft_SDFChainRadix22__T_400) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_411 = fft_fft_SDFChainRadix22__T_410[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_418 = fft_fft_SDFChainRadix22_sdf_stages_4_io_cntr < 9'h10; // @[SDFChainRadix22.scala 328:32]
  assign fft_fft_SDFChainRadix22__T_419 = fft_fft_SDFChainRadix22_sdf_stages_4_io_cntr < 9'h18; // @[SDFChainRadix22.scala 328:78]
  assign fft_fft_SDFChainRadix22__T_420 = fft_fft_SDFChainRadix22__T_419 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign fft_fft_SDFChainRadix22__T_421 = fft_fft_SDFChainRadix22__T_418 ? 1'h0 : fft_fft_SDFChainRadix22__T_420; // @[SDFChainRadix22.scala 328:19]
  assign fft_fft_SDFChainRadix22_outputWires_3_real = fft_fft_SDFChainRadix22_sdf_stages_3_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__T_427 = 16'sh0 - $signed(fft_fft_SDFChainRadix22_outputWires_3_real); // @[FixedPointTypeClass.scala 39:43]
  assign fft_fft_SDFChainRadix22_outputWires_3_imag = fft_fft_SDFChainRadix22_sdf_stages_3_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__T_759 = fft_fft_SDFChainRadix22__T_201[6:0];
  assign fft_fft_SDFChainRadix22__GEN_202 = 7'h21 == fft_fft_SDFChainRadix22__T_759 ? 6'h2 : 6'h0; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_203 = 7'h22 == fft_fft_SDFChainRadix22__T_759 ? 6'h4 : fft_fft_SDFChainRadix22__GEN_202; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_204 = 7'h23 == fft_fft_SDFChainRadix22__T_759 ? 6'h6 : fft_fft_SDFChainRadix22__GEN_203; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_205 = 7'h24 == fft_fft_SDFChainRadix22__T_759 ? 6'h8 : fft_fft_SDFChainRadix22__GEN_204; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_206 = 7'h25 == fft_fft_SDFChainRadix22__T_759 ? 6'ha : fft_fft_SDFChainRadix22__GEN_205; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_207 = 7'h26 == fft_fft_SDFChainRadix22__T_759 ? 6'hc : fft_fft_SDFChainRadix22__GEN_206; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_208 = 7'h27 == fft_fft_SDFChainRadix22__T_759 ? 6'he : fft_fft_SDFChainRadix22__GEN_207; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_209 = 7'h28 == fft_fft_SDFChainRadix22__T_759 ? 6'h10 : fft_fft_SDFChainRadix22__GEN_208; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_210 = 7'h29 == fft_fft_SDFChainRadix22__T_759 ? 6'h12 : fft_fft_SDFChainRadix22__GEN_209; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_211 = 7'h2a == fft_fft_SDFChainRadix22__T_759 ? 6'h14 : fft_fft_SDFChainRadix22__GEN_210; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_212 = 7'h2b == fft_fft_SDFChainRadix22__T_759 ? 6'h16 : fft_fft_SDFChainRadix22__GEN_211; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_213 = 7'h2c == fft_fft_SDFChainRadix22__T_759 ? 6'h18 : fft_fft_SDFChainRadix22__GEN_212; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_214 = 7'h2d == fft_fft_SDFChainRadix22__T_759 ? 6'h1a : fft_fft_SDFChainRadix22__GEN_213; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_215 = 7'h2e == fft_fft_SDFChainRadix22__T_759 ? 6'h1c : fft_fft_SDFChainRadix22__GEN_214; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_216 = 7'h2f == fft_fft_SDFChainRadix22__T_759 ? 6'h1e : fft_fft_SDFChainRadix22__GEN_215; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_217 = 7'h30 == fft_fft_SDFChainRadix22__T_759 ? 6'h20 : fft_fft_SDFChainRadix22__GEN_216; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_218 = 7'h31 == fft_fft_SDFChainRadix22__T_759 ? 6'h22 : fft_fft_SDFChainRadix22__GEN_217; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_219 = 7'h32 == fft_fft_SDFChainRadix22__T_759 ? 6'h23 : fft_fft_SDFChainRadix22__GEN_218; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_220 = 7'h33 == fft_fft_SDFChainRadix22__T_759 ? 6'h24 : fft_fft_SDFChainRadix22__GEN_219; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_221 = 7'h34 == fft_fft_SDFChainRadix22__T_759 ? 6'h26 : fft_fft_SDFChainRadix22__GEN_220; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_222 = 7'h35 == fft_fft_SDFChainRadix22__T_759 ? 6'h27 : fft_fft_SDFChainRadix22__GEN_221; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_223 = 7'h36 == fft_fft_SDFChainRadix22__T_759 ? 6'h28 : fft_fft_SDFChainRadix22__GEN_222; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_224 = 7'h37 == fft_fft_SDFChainRadix22__T_759 ? 6'h2a : fft_fft_SDFChainRadix22__GEN_223; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_225 = 7'h38 == fft_fft_SDFChainRadix22__T_759 ? 6'h2b : fft_fft_SDFChainRadix22__GEN_224; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_226 = 7'h39 == fft_fft_SDFChainRadix22__T_759 ? 6'h2c : fft_fft_SDFChainRadix22__GEN_225; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_227 = 7'h3a == fft_fft_SDFChainRadix22__T_759 ? 6'h2e : fft_fft_SDFChainRadix22__GEN_226; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_228 = 7'h3b == fft_fft_SDFChainRadix22__T_759 ? 6'h2f : fft_fft_SDFChainRadix22__GEN_227; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_229 = 7'h3c == fft_fft_SDFChainRadix22__T_759 ? 6'h30 : fft_fft_SDFChainRadix22__GEN_228; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_230 = 7'h3d == fft_fft_SDFChainRadix22__T_759 ? 6'h32 : fft_fft_SDFChainRadix22__GEN_229; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_231 = 7'h3e == fft_fft_SDFChainRadix22__T_759 ? 6'h33 : fft_fft_SDFChainRadix22__GEN_230; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_232 = 7'h3f == fft_fft_SDFChainRadix22__T_759 ? 6'h34 : fft_fft_SDFChainRadix22__GEN_231; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_233 = 7'h40 == fft_fft_SDFChainRadix22__T_759 ? 6'h0 : fft_fft_SDFChainRadix22__GEN_232; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_234 = 7'h41 == fft_fft_SDFChainRadix22__T_759 ? 6'h1 : fft_fft_SDFChainRadix22__GEN_233; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_235 = 7'h42 == fft_fft_SDFChainRadix22__T_759 ? 6'h2 : fft_fft_SDFChainRadix22__GEN_234; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_236 = 7'h43 == fft_fft_SDFChainRadix22__T_759 ? 6'h3 : fft_fft_SDFChainRadix22__GEN_235; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_237 = 7'h44 == fft_fft_SDFChainRadix22__T_759 ? 6'h4 : fft_fft_SDFChainRadix22__GEN_236; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_238 = 7'h45 == fft_fft_SDFChainRadix22__T_759 ? 6'h5 : fft_fft_SDFChainRadix22__GEN_237; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_239 = 7'h46 == fft_fft_SDFChainRadix22__T_759 ? 6'h6 : fft_fft_SDFChainRadix22__GEN_238; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_240 = 7'h47 == fft_fft_SDFChainRadix22__T_759 ? 6'h7 : fft_fft_SDFChainRadix22__GEN_239; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_241 = 7'h48 == fft_fft_SDFChainRadix22__T_759 ? 6'h8 : fft_fft_SDFChainRadix22__GEN_240; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_242 = 7'h49 == fft_fft_SDFChainRadix22__T_759 ? 6'h9 : fft_fft_SDFChainRadix22__GEN_241; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_243 = 7'h4a == fft_fft_SDFChainRadix22__T_759 ? 6'ha : fft_fft_SDFChainRadix22__GEN_242; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_244 = 7'h4b == fft_fft_SDFChainRadix22__T_759 ? 6'hb : fft_fft_SDFChainRadix22__GEN_243; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_245 = 7'h4c == fft_fft_SDFChainRadix22__T_759 ? 6'hc : fft_fft_SDFChainRadix22__GEN_244; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_246 = 7'h4d == fft_fft_SDFChainRadix22__T_759 ? 6'hd : fft_fft_SDFChainRadix22__GEN_245; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_247 = 7'h4e == fft_fft_SDFChainRadix22__T_759 ? 6'he : fft_fft_SDFChainRadix22__GEN_246; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_248 = 7'h4f == fft_fft_SDFChainRadix22__T_759 ? 6'hf : fft_fft_SDFChainRadix22__GEN_247; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_249 = 7'h50 == fft_fft_SDFChainRadix22__T_759 ? 6'h10 : fft_fft_SDFChainRadix22__GEN_248; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_250 = 7'h51 == fft_fft_SDFChainRadix22__T_759 ? 6'h11 : fft_fft_SDFChainRadix22__GEN_249; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_251 = 7'h52 == fft_fft_SDFChainRadix22__T_759 ? 6'h12 : fft_fft_SDFChainRadix22__GEN_250; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_252 = 7'h53 == fft_fft_SDFChainRadix22__T_759 ? 6'h13 : fft_fft_SDFChainRadix22__GEN_251; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_253 = 7'h54 == fft_fft_SDFChainRadix22__T_759 ? 6'h14 : fft_fft_SDFChainRadix22__GEN_252; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_254 = 7'h55 == fft_fft_SDFChainRadix22__T_759 ? 6'h15 : fft_fft_SDFChainRadix22__GEN_253; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_255 = 7'h56 == fft_fft_SDFChainRadix22__T_759 ? 6'h16 : fft_fft_SDFChainRadix22__GEN_254; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_256 = 7'h57 == fft_fft_SDFChainRadix22__T_759 ? 6'h17 : fft_fft_SDFChainRadix22__GEN_255; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_257 = 7'h58 == fft_fft_SDFChainRadix22__T_759 ? 6'h18 : fft_fft_SDFChainRadix22__GEN_256; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_258 = 7'h59 == fft_fft_SDFChainRadix22__T_759 ? 6'h19 : fft_fft_SDFChainRadix22__GEN_257; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_259 = 7'h5a == fft_fft_SDFChainRadix22__T_759 ? 6'h1a : fft_fft_SDFChainRadix22__GEN_258; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_260 = 7'h5b == fft_fft_SDFChainRadix22__T_759 ? 6'h1b : fft_fft_SDFChainRadix22__GEN_259; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_261 = 7'h5c == fft_fft_SDFChainRadix22__T_759 ? 6'h1c : fft_fft_SDFChainRadix22__GEN_260; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_262 = 7'h5d == fft_fft_SDFChainRadix22__T_759 ? 6'h1d : fft_fft_SDFChainRadix22__GEN_261; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_263 = 7'h5e == fft_fft_SDFChainRadix22__T_759 ? 6'h1e : fft_fft_SDFChainRadix22__GEN_262; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_264 = 7'h5f == fft_fft_SDFChainRadix22__T_759 ? 6'h1f : fft_fft_SDFChainRadix22__GEN_263; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_265 = 7'h60 == fft_fft_SDFChainRadix22__T_759 ? 6'h0 : fft_fft_SDFChainRadix22__GEN_264; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_266 = 7'h61 == fft_fft_SDFChainRadix22__T_759 ? 6'h3 : fft_fft_SDFChainRadix22__GEN_265; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_267 = 7'h62 == fft_fft_SDFChainRadix22__T_759 ? 6'h6 : fft_fft_SDFChainRadix22__GEN_266; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_268 = 7'h63 == fft_fft_SDFChainRadix22__T_759 ? 6'h9 : fft_fft_SDFChainRadix22__GEN_267; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_269 = 7'h64 == fft_fft_SDFChainRadix22__T_759 ? 6'hc : fft_fft_SDFChainRadix22__GEN_268; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_270 = 7'h65 == fft_fft_SDFChainRadix22__T_759 ? 6'hf : fft_fft_SDFChainRadix22__GEN_269; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_271 = 7'h66 == fft_fft_SDFChainRadix22__T_759 ? 6'h12 : fft_fft_SDFChainRadix22__GEN_270; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_272 = 7'h67 == fft_fft_SDFChainRadix22__T_759 ? 6'h15 : fft_fft_SDFChainRadix22__GEN_271; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_273 = 7'h68 == fft_fft_SDFChainRadix22__T_759 ? 6'h18 : fft_fft_SDFChainRadix22__GEN_272; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_274 = 7'h69 == fft_fft_SDFChainRadix22__T_759 ? 6'h1b : fft_fft_SDFChainRadix22__GEN_273; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_275 = 7'h6a == fft_fft_SDFChainRadix22__T_759 ? 6'h1e : fft_fft_SDFChainRadix22__GEN_274; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_276 = 7'h6b == fft_fft_SDFChainRadix22__T_759 ? 6'h21 : fft_fft_SDFChainRadix22__GEN_275; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_277 = 7'h6c == fft_fft_SDFChainRadix22__T_759 ? 6'h23 : fft_fft_SDFChainRadix22__GEN_276; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_278 = 7'h6d == fft_fft_SDFChainRadix22__T_759 ? 6'h25 : fft_fft_SDFChainRadix22__GEN_277; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_279 = 7'h6e == fft_fft_SDFChainRadix22__T_759 ? 6'h27 : fft_fft_SDFChainRadix22__GEN_278; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_280 = 7'h6f == fft_fft_SDFChainRadix22__T_759 ? 6'h29 : fft_fft_SDFChainRadix22__GEN_279; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_281 = 7'h70 == fft_fft_SDFChainRadix22__T_759 ? 6'h2b : fft_fft_SDFChainRadix22__GEN_280; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_282 = 7'h71 == fft_fft_SDFChainRadix22__T_759 ? 6'h2d : fft_fft_SDFChainRadix22__GEN_281; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_283 = 7'h72 == fft_fft_SDFChainRadix22__T_759 ? 6'h2f : fft_fft_SDFChainRadix22__GEN_282; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_284 = 7'h73 == fft_fft_SDFChainRadix22__T_759 ? 6'h31 : fft_fft_SDFChainRadix22__GEN_283; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_285 = 7'h74 == fft_fft_SDFChainRadix22__T_759 ? 6'h33 : fft_fft_SDFChainRadix22__GEN_284; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_286 = 7'h75 == fft_fft_SDFChainRadix22__T_759 ? 6'h35 : fft_fft_SDFChainRadix22__GEN_285; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_287 = 7'h76 == fft_fft_SDFChainRadix22__T_759 ? 6'h36 : fft_fft_SDFChainRadix22__GEN_286; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_288 = 7'h77 == fft_fft_SDFChainRadix22__T_759 ? 6'h37 : fft_fft_SDFChainRadix22__GEN_287; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_289 = 7'h78 == fft_fft_SDFChainRadix22__T_759 ? 6'h38 : fft_fft_SDFChainRadix22__GEN_288; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_290 = 7'h79 == fft_fft_SDFChainRadix22__T_759 ? 6'h39 : fft_fft_SDFChainRadix22__GEN_289; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_291 = 7'h7a == fft_fft_SDFChainRadix22__T_759 ? 6'h3a : fft_fft_SDFChainRadix22__GEN_290; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_292 = 7'h7b == fft_fft_SDFChainRadix22__T_759 ? 6'h3b : fft_fft_SDFChainRadix22__GEN_291; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_293 = 7'h7c == fft_fft_SDFChainRadix22__T_759 ? 6'h3c : fft_fft_SDFChainRadix22__GEN_292; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_294 = 7'h7d == fft_fft_SDFChainRadix22__T_759 ? 6'h3d : fft_fft_SDFChainRadix22__GEN_293; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_295 = 7'h7e == fft_fft_SDFChainRadix22__T_759 ? 6'h3e : fft_fft_SDFChainRadix22__GEN_294; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_296 = 7'h7f == fft_fft_SDFChainRadix22__T_759 ? 6'h3f : fft_fft_SDFChainRadix22__GEN_295; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_299 = 6'h1 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3fec) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_300 = 6'h1 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh324) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_301 = 6'h2 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_299); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_302 = 6'h2 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_300); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_303 = 6'h3 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_301); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_304 = 6'h3 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_302); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_305 = 6'h4 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_303); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_306 = 6'h4 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_304); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_307 = 6'h5 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_305); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_308 = 6'h5 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_306); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_309 = 6'h6 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_307); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_310 = 6'h6 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_308); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_311 = 6'h7 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_309); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_312 = 6'h7 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_310); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_313 = 6'h8 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_311); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_314 = 6'h8 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_312); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_315 = 6'h9 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_313); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_316 = 6'h9 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_314); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_317 = 6'ha == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_315); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_318 = 6'ha == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_316); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_319 = 6'hb == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_317); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_320 = 6'hb == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_318); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_321 = 6'hc == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_319); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_322 = 6'hc == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_320); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_323 = 6'hd == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_321); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_324 = 6'hd == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_322); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_325 = 6'he == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_323); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_326 = 6'he == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_324); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_327 = 6'hf == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_325); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_328 = 6'hf == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_326); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_329 = 6'h10 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_327); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_330 = 6'h10 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_328); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_331 = 6'h11 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_329); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_332 = 6'h11 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_330); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_333 = 6'h12 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_331); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_334 = 6'h12 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_332); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_335 = 6'h13 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_333); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_336 = 6'h13 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_334); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_337 = 6'h14 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_335); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_338 = 6'h14 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_336); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_339 = 6'h15 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_337); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_340 = 6'h15 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_338); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_341 = 6'h16 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_339); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_342 = 6'h16 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_340); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_343 = 6'h17 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_341); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_344 = 6'h17 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_342); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_345 = 6'h18 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_343); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_346 = 6'h18 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_344); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_347 = 6'h19 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_345); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_348 = 6'h19 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_346); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_349 = 6'h1a == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_347); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_350 = 6'h1a == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_348); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_351 = 6'h1b == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_349); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_352 = 6'h1b == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_350); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_353 = 6'h1c == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_351); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_354 = 6'h1c == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_352); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_355 = 6'h1d == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_353); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_356 = 6'h1d == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_354); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_357 = 6'h1e == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_355); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_358 = 6'h1e == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_356); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_359 = 6'h1f == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh324) : $signed(fft_fft_SDFChainRadix22__GEN_357); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_360 = 6'h1f == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3fec) : $signed(fft_fft_SDFChainRadix22__GEN_358); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_361 = 6'h20 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh0) : $signed(fft_fft_SDFChainRadix22__GEN_359); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_362 = 6'h20 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh4000) : $signed(fft_fft_SDFChainRadix22__GEN_360); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_363 = 6'h21 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh324) : $signed(fft_fft_SDFChainRadix22__GEN_361); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_364 = 6'h21 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3fec) : $signed(fft_fft_SDFChainRadix22__GEN_362); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_365 = 6'h22 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_363); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_366 = 6'h22 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_364); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_367 = 6'h23 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_365); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_368 = 6'h23 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_366); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_369 = 6'h24 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_367); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_370 = 6'h24 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_368); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_371 = 6'h25 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_369); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_372 = 6'h25 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_370); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_373 = 6'h26 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_371); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_374 = 6'h26 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_372); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_375 = 6'h27 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_373); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_376 = 6'h27 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_374); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_377 = 6'h28 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_375); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_378 = 6'h28 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_376); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_379 = 6'h29 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_377); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_380 = 6'h29 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_378); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_381 = 6'h2a == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_379); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_382 = 6'h2a == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_380); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_383 = 6'h2b == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_381); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_384 = 6'h2b == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_382); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_385 = 6'h2c == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_383); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_386 = 6'h2c == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_384); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_387 = 6'h2d == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_385); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_388 = 6'h2d == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_386); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_389 = 6'h2e == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_387); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_390 = 6'h2e == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_388); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_391 = 6'h2f == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_389); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_392 = 6'h2f == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_390); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_393 = 6'h30 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_391); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_394 = 6'h30 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_392); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_395 = 6'h31 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_393); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_396 = 6'h31 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_394); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_397 = 6'h32 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_395); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_398 = 6'h32 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_396); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_399 = 6'h33 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_397); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_400 = 6'h33 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_398); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_401 = 6'h34 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_399); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_402 = 6'h34 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_400); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_403 = 6'h35 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3fec) : $signed(fft_fft_SDFChainRadix22__GEN_401); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_404 = 6'h35 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh324) : $signed(fft_fft_SDFChainRadix22__GEN_402); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_405 = 6'h36 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_403); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_406 = 6'h36 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_404); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_407 = 6'h37 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_405); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_408 = 6'h37 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_406); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_409 = 6'h38 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_407); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_410 = 6'h38 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_408); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_411 = 6'h39 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_409); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_412 = 6'h39 == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_410); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_413 = 6'h3a == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_411); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_414 = 6'h3a == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_412); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_415 = 6'h3b == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_413); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_416 = 6'h3b == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_414); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_417 = 6'h3c == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_415); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_418 = 6'h3c == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_416); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_419 = 6'h3d == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_417); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_420 = 6'h3d == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_418); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_421 = 6'h3e == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_419); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_422 = 6'h3e == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_420); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_423 = 6'h3f == fft_fft_SDFChainRadix22__GEN_296 ? $signed(-16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_421); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22_twiddles_5_imag = 6'h3f == fft_fft_SDFChainRadix22__GEN_296 ? $signed(16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_422); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__T_765 = $signed(fft_fft_SDFChainRadix22__GEN_423) + $signed(fft_fft_SDFChainRadix22_twiddles_5_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_outputWires_4_real = fft_fft_SDFChainRadix22_sdf_stages_4_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22_outputWires_4_imag = fft_fft_SDFChainRadix22_sdf_stages_4_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22__T_766 = $signed(fft_fft_SDFChainRadix22_outputWires_4_real) + $signed(fft_fft_SDFChainRadix22_outputWires_4_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_767 = $signed(fft_fft_SDFChainRadix22_outputWires_4_imag) - $signed(fft_fft_SDFChainRadix22_outputWires_4_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__GEN_2118 = {{1{fft_fft_SDFChainRadix22_outputWires_4_real[15]}},fft_fft_SDFChainRadix22_outputWires_4_real}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_768 = $signed(fft_fft_SDFChainRadix22__GEN_2118) * $signed(fft_fft_SDFChainRadix22__T_765); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2119 = {{1{fft_fft_SDFChainRadix22_twiddles_5_imag[15]}},fft_fft_SDFChainRadix22_twiddles_5_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_769 = $signed(fft_fft_SDFChainRadix22__T_766) * $signed(fft_fft_SDFChainRadix22__GEN_2119); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2120 = {{1{fft_fft_SDFChainRadix22__GEN_423[15]}},fft_fft_SDFChainRadix22__GEN_423}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_770 = $signed(fft_fft_SDFChainRadix22__T_767) * $signed(fft_fft_SDFChainRadix22__GEN_2120); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_771 = $signed(fft_fft_SDFChainRadix22__T_768) - $signed(fft_fft_SDFChainRadix22__T_769); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__T_772 = $signed(fft_fft_SDFChainRadix22__T_768) + $signed(fft_fft_SDFChainRadix22__T_770); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_778 = $signed(fft_fft_SDFChainRadix22__T_771) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_779 = fft_fft_SDFChainRadix22__T_778[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_782 = $signed(fft_fft_SDFChainRadix22__T_772) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_783 = fft_fft_SDFChainRadix22__T_782[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_790 = fft_fft_SDFChainRadix22_sdf_stages_6_io_cntr < 9'h40; // @[SDFChainRadix22.scala 328:32]
  assign fft_fft_SDFChainRadix22__T_791 = fft_fft_SDFChainRadix22_sdf_stages_6_io_cntr < 9'h60; // @[SDFChainRadix22.scala 328:78]
  assign fft_fft_SDFChainRadix22__T_792 = fft_fft_SDFChainRadix22__T_791 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign fft_fft_SDFChainRadix22__T_793 = fft_fft_SDFChainRadix22__T_790 ? 1'h0 : fft_fft_SDFChainRadix22__T_792; // @[SDFChainRadix22.scala 328:19]
  assign fft_fft_SDFChainRadix22_outputWires_5_real = fft_fft_SDFChainRadix22_sdf_stages_5_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__T_799 = 16'sh0 - $signed(fft_fft_SDFChainRadix22_outputWires_5_real); // @[FixedPointTypeClass.scala 39:43]
  assign fft_fft_SDFChainRadix22_outputWires_5_imag = fft_fft_SDFChainRadix22_sdf_stages_5_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__GEN_682 = 9'h81 == fft_fft_SDFChainRadix22__T_215 ? 8'h2 : 8'h0; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_683 = 9'h82 == fft_fft_SDFChainRadix22__T_215 ? 8'h4 : fft_fft_SDFChainRadix22__GEN_682; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_684 = 9'h83 == fft_fft_SDFChainRadix22__T_215 ? 8'h6 : fft_fft_SDFChainRadix22__GEN_683; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_685 = 9'h84 == fft_fft_SDFChainRadix22__T_215 ? 8'h8 : fft_fft_SDFChainRadix22__GEN_684; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_686 = 9'h85 == fft_fft_SDFChainRadix22__T_215 ? 8'ha : fft_fft_SDFChainRadix22__GEN_685; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_687 = 9'h86 == fft_fft_SDFChainRadix22__T_215 ? 8'hc : fft_fft_SDFChainRadix22__GEN_686; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_688 = 9'h87 == fft_fft_SDFChainRadix22__T_215 ? 8'he : fft_fft_SDFChainRadix22__GEN_687; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_689 = 9'h88 == fft_fft_SDFChainRadix22__T_215 ? 8'h10 : fft_fft_SDFChainRadix22__GEN_688; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_690 = 9'h89 == fft_fft_SDFChainRadix22__T_215 ? 8'h12 : fft_fft_SDFChainRadix22__GEN_689; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_691 = 9'h8a == fft_fft_SDFChainRadix22__T_215 ? 8'h14 : fft_fft_SDFChainRadix22__GEN_690; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_692 = 9'h8b == fft_fft_SDFChainRadix22__T_215 ? 8'h16 : fft_fft_SDFChainRadix22__GEN_691; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_693 = 9'h8c == fft_fft_SDFChainRadix22__T_215 ? 8'h18 : fft_fft_SDFChainRadix22__GEN_692; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_694 = 9'h8d == fft_fft_SDFChainRadix22__T_215 ? 8'h1a : fft_fft_SDFChainRadix22__GEN_693; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_695 = 9'h8e == fft_fft_SDFChainRadix22__T_215 ? 8'h1c : fft_fft_SDFChainRadix22__GEN_694; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_696 = 9'h8f == fft_fft_SDFChainRadix22__T_215 ? 8'h1e : fft_fft_SDFChainRadix22__GEN_695; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_697 = 9'h90 == fft_fft_SDFChainRadix22__T_215 ? 8'h20 : fft_fft_SDFChainRadix22__GEN_696; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_698 = 9'h91 == fft_fft_SDFChainRadix22__T_215 ? 8'h22 : fft_fft_SDFChainRadix22__GEN_697; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_699 = 9'h92 == fft_fft_SDFChainRadix22__T_215 ? 8'h24 : fft_fft_SDFChainRadix22__GEN_698; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_700 = 9'h93 == fft_fft_SDFChainRadix22__T_215 ? 8'h26 : fft_fft_SDFChainRadix22__GEN_699; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_701 = 9'h94 == fft_fft_SDFChainRadix22__T_215 ? 8'h28 : fft_fft_SDFChainRadix22__GEN_700; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_702 = 9'h95 == fft_fft_SDFChainRadix22__T_215 ? 8'h2a : fft_fft_SDFChainRadix22__GEN_701; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_703 = 9'h96 == fft_fft_SDFChainRadix22__T_215 ? 8'h2c : fft_fft_SDFChainRadix22__GEN_702; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_704 = 9'h97 == fft_fft_SDFChainRadix22__T_215 ? 8'h2e : fft_fft_SDFChainRadix22__GEN_703; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_705 = 9'h98 == fft_fft_SDFChainRadix22__T_215 ? 8'h30 : fft_fft_SDFChainRadix22__GEN_704; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_706 = 9'h99 == fft_fft_SDFChainRadix22__T_215 ? 8'h32 : fft_fft_SDFChainRadix22__GEN_705; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_707 = 9'h9a == fft_fft_SDFChainRadix22__T_215 ? 8'h34 : fft_fft_SDFChainRadix22__GEN_706; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_708 = 9'h9b == fft_fft_SDFChainRadix22__T_215 ? 8'h36 : fft_fft_SDFChainRadix22__GEN_707; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_709 = 9'h9c == fft_fft_SDFChainRadix22__T_215 ? 8'h38 : fft_fft_SDFChainRadix22__GEN_708; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_710 = 9'h9d == fft_fft_SDFChainRadix22__T_215 ? 8'h3a : fft_fft_SDFChainRadix22__GEN_709; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_711 = 9'h9e == fft_fft_SDFChainRadix22__T_215 ? 8'h3c : fft_fft_SDFChainRadix22__GEN_710; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_712 = 9'h9f == fft_fft_SDFChainRadix22__T_215 ? 8'h3e : fft_fft_SDFChainRadix22__GEN_711; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_713 = 9'ha0 == fft_fft_SDFChainRadix22__T_215 ? 8'h40 : fft_fft_SDFChainRadix22__GEN_712; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_714 = 9'ha1 == fft_fft_SDFChainRadix22__T_215 ? 8'h42 : fft_fft_SDFChainRadix22__GEN_713; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_715 = 9'ha2 == fft_fft_SDFChainRadix22__T_215 ? 8'h44 : fft_fft_SDFChainRadix22__GEN_714; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_716 = 9'ha3 == fft_fft_SDFChainRadix22__T_215 ? 8'h46 : fft_fft_SDFChainRadix22__GEN_715; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_717 = 9'ha4 == fft_fft_SDFChainRadix22__T_215 ? 8'h48 : fft_fft_SDFChainRadix22__GEN_716; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_718 = 9'ha5 == fft_fft_SDFChainRadix22__T_215 ? 8'h4a : fft_fft_SDFChainRadix22__GEN_717; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_719 = 9'ha6 == fft_fft_SDFChainRadix22__T_215 ? 8'h4c : fft_fft_SDFChainRadix22__GEN_718; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_720 = 9'ha7 == fft_fft_SDFChainRadix22__T_215 ? 8'h4e : fft_fft_SDFChainRadix22__GEN_719; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_721 = 9'ha8 == fft_fft_SDFChainRadix22__T_215 ? 8'h50 : fft_fft_SDFChainRadix22__GEN_720; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_722 = 9'ha9 == fft_fft_SDFChainRadix22__T_215 ? 8'h52 : fft_fft_SDFChainRadix22__GEN_721; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_723 = 9'haa == fft_fft_SDFChainRadix22__T_215 ? 8'h54 : fft_fft_SDFChainRadix22__GEN_722; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_724 = 9'hab == fft_fft_SDFChainRadix22__T_215 ? 8'h56 : fft_fft_SDFChainRadix22__GEN_723; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_725 = 9'hac == fft_fft_SDFChainRadix22__T_215 ? 8'h58 : fft_fft_SDFChainRadix22__GEN_724; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_726 = 9'had == fft_fft_SDFChainRadix22__T_215 ? 8'h5a : fft_fft_SDFChainRadix22__GEN_725; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_727 = 9'hae == fft_fft_SDFChainRadix22__T_215 ? 8'h5c : fft_fft_SDFChainRadix22__GEN_726; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_728 = 9'haf == fft_fft_SDFChainRadix22__T_215 ? 8'h5e : fft_fft_SDFChainRadix22__GEN_727; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_729 = 9'hb0 == fft_fft_SDFChainRadix22__T_215 ? 8'h60 : fft_fft_SDFChainRadix22__GEN_728; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_730 = 9'hb1 == fft_fft_SDFChainRadix22__T_215 ? 8'h62 : fft_fft_SDFChainRadix22__GEN_729; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_731 = 9'hb2 == fft_fft_SDFChainRadix22__T_215 ? 8'h64 : fft_fft_SDFChainRadix22__GEN_730; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_732 = 9'hb3 == fft_fft_SDFChainRadix22__T_215 ? 8'h66 : fft_fft_SDFChainRadix22__GEN_731; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_733 = 9'hb4 == fft_fft_SDFChainRadix22__T_215 ? 8'h68 : fft_fft_SDFChainRadix22__GEN_732; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_734 = 9'hb5 == fft_fft_SDFChainRadix22__T_215 ? 8'h6a : fft_fft_SDFChainRadix22__GEN_733; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_735 = 9'hb6 == fft_fft_SDFChainRadix22__T_215 ? 8'h6c : fft_fft_SDFChainRadix22__GEN_734; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_736 = 9'hb7 == fft_fft_SDFChainRadix22__T_215 ? 8'h6e : fft_fft_SDFChainRadix22__GEN_735; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_737 = 9'hb8 == fft_fft_SDFChainRadix22__T_215 ? 8'h70 : fft_fft_SDFChainRadix22__GEN_736; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_738 = 9'hb9 == fft_fft_SDFChainRadix22__T_215 ? 8'h72 : fft_fft_SDFChainRadix22__GEN_737; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_739 = 9'hba == fft_fft_SDFChainRadix22__T_215 ? 8'h74 : fft_fft_SDFChainRadix22__GEN_738; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_740 = 9'hbb == fft_fft_SDFChainRadix22__T_215 ? 8'h76 : fft_fft_SDFChainRadix22__GEN_739; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_741 = 9'hbc == fft_fft_SDFChainRadix22__T_215 ? 8'h78 : fft_fft_SDFChainRadix22__GEN_740; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_742 = 9'hbd == fft_fft_SDFChainRadix22__T_215 ? 8'h7a : fft_fft_SDFChainRadix22__GEN_741; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_743 = 9'hbe == fft_fft_SDFChainRadix22__T_215 ? 8'h7c : fft_fft_SDFChainRadix22__GEN_742; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_744 = 9'hbf == fft_fft_SDFChainRadix22__T_215 ? 8'h7e : fft_fft_SDFChainRadix22__GEN_743; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_745 = 9'hc0 == fft_fft_SDFChainRadix22__T_215 ? 8'h80 : fft_fft_SDFChainRadix22__GEN_744; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_746 = 9'hc1 == fft_fft_SDFChainRadix22__T_215 ? 8'h82 : fft_fft_SDFChainRadix22__GEN_745; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_747 = 9'hc2 == fft_fft_SDFChainRadix22__T_215 ? 8'h83 : fft_fft_SDFChainRadix22__GEN_746; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_748 = 9'hc3 == fft_fft_SDFChainRadix22__T_215 ? 8'h84 : fft_fft_SDFChainRadix22__GEN_747; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_749 = 9'hc4 == fft_fft_SDFChainRadix22__T_215 ? 8'h86 : fft_fft_SDFChainRadix22__GEN_748; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_750 = 9'hc5 == fft_fft_SDFChainRadix22__T_215 ? 8'h87 : fft_fft_SDFChainRadix22__GEN_749; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_751 = 9'hc6 == fft_fft_SDFChainRadix22__T_215 ? 8'h88 : fft_fft_SDFChainRadix22__GEN_750; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_752 = 9'hc7 == fft_fft_SDFChainRadix22__T_215 ? 8'h8a : fft_fft_SDFChainRadix22__GEN_751; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_753 = 9'hc8 == fft_fft_SDFChainRadix22__T_215 ? 8'h8b : fft_fft_SDFChainRadix22__GEN_752; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_754 = 9'hc9 == fft_fft_SDFChainRadix22__T_215 ? 8'h8c : fft_fft_SDFChainRadix22__GEN_753; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_755 = 9'hca == fft_fft_SDFChainRadix22__T_215 ? 8'h8e : fft_fft_SDFChainRadix22__GEN_754; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_756 = 9'hcb == fft_fft_SDFChainRadix22__T_215 ? 8'h8f : fft_fft_SDFChainRadix22__GEN_755; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_757 = 9'hcc == fft_fft_SDFChainRadix22__T_215 ? 8'h90 : fft_fft_SDFChainRadix22__GEN_756; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_758 = 9'hcd == fft_fft_SDFChainRadix22__T_215 ? 8'h92 : fft_fft_SDFChainRadix22__GEN_757; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_759 = 9'hce == fft_fft_SDFChainRadix22__T_215 ? 8'h93 : fft_fft_SDFChainRadix22__GEN_758; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_760 = 9'hcf == fft_fft_SDFChainRadix22__T_215 ? 8'h94 : fft_fft_SDFChainRadix22__GEN_759; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_761 = 9'hd0 == fft_fft_SDFChainRadix22__T_215 ? 8'h96 : fft_fft_SDFChainRadix22__GEN_760; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_762 = 9'hd1 == fft_fft_SDFChainRadix22__T_215 ? 8'h97 : fft_fft_SDFChainRadix22__GEN_761; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_763 = 9'hd2 == fft_fft_SDFChainRadix22__T_215 ? 8'h98 : fft_fft_SDFChainRadix22__GEN_762; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_764 = 9'hd3 == fft_fft_SDFChainRadix22__T_215 ? 8'h9a : fft_fft_SDFChainRadix22__GEN_763; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_765 = 9'hd4 == fft_fft_SDFChainRadix22__T_215 ? 8'h9b : fft_fft_SDFChainRadix22__GEN_764; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_766 = 9'hd5 == fft_fft_SDFChainRadix22__T_215 ? 8'h9c : fft_fft_SDFChainRadix22__GEN_765; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_767 = 9'hd6 == fft_fft_SDFChainRadix22__T_215 ? 8'h9e : fft_fft_SDFChainRadix22__GEN_766; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_768 = 9'hd7 == fft_fft_SDFChainRadix22__T_215 ? 8'h9f : fft_fft_SDFChainRadix22__GEN_767; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_769 = 9'hd8 == fft_fft_SDFChainRadix22__T_215 ? 8'ha0 : fft_fft_SDFChainRadix22__GEN_768; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_770 = 9'hd9 == fft_fft_SDFChainRadix22__T_215 ? 8'ha2 : fft_fft_SDFChainRadix22__GEN_769; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_771 = 9'hda == fft_fft_SDFChainRadix22__T_215 ? 8'ha3 : fft_fft_SDFChainRadix22__GEN_770; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_772 = 9'hdb == fft_fft_SDFChainRadix22__T_215 ? 8'ha4 : fft_fft_SDFChainRadix22__GEN_771; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_773 = 9'hdc == fft_fft_SDFChainRadix22__T_215 ? 8'ha6 : fft_fft_SDFChainRadix22__GEN_772; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_774 = 9'hdd == fft_fft_SDFChainRadix22__T_215 ? 8'ha7 : fft_fft_SDFChainRadix22__GEN_773; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_775 = 9'hde == fft_fft_SDFChainRadix22__T_215 ? 8'ha8 : fft_fft_SDFChainRadix22__GEN_774; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_776 = 9'hdf == fft_fft_SDFChainRadix22__T_215 ? 8'haa : fft_fft_SDFChainRadix22__GEN_775; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_777 = 9'he0 == fft_fft_SDFChainRadix22__T_215 ? 8'hab : fft_fft_SDFChainRadix22__GEN_776; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_778 = 9'he1 == fft_fft_SDFChainRadix22__T_215 ? 8'hac : fft_fft_SDFChainRadix22__GEN_777; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_779 = 9'he2 == fft_fft_SDFChainRadix22__T_215 ? 8'hae : fft_fft_SDFChainRadix22__GEN_778; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_780 = 9'he3 == fft_fft_SDFChainRadix22__T_215 ? 8'haf : fft_fft_SDFChainRadix22__GEN_779; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_781 = 9'he4 == fft_fft_SDFChainRadix22__T_215 ? 8'hb0 : fft_fft_SDFChainRadix22__GEN_780; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_782 = 9'he5 == fft_fft_SDFChainRadix22__T_215 ? 8'hb2 : fft_fft_SDFChainRadix22__GEN_781; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_783 = 9'he6 == fft_fft_SDFChainRadix22__T_215 ? 8'hb3 : fft_fft_SDFChainRadix22__GEN_782; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_784 = 9'he7 == fft_fft_SDFChainRadix22__T_215 ? 8'hb4 : fft_fft_SDFChainRadix22__GEN_783; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_785 = 9'he8 == fft_fft_SDFChainRadix22__T_215 ? 8'hb6 : fft_fft_SDFChainRadix22__GEN_784; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_786 = 9'he9 == fft_fft_SDFChainRadix22__T_215 ? 8'hb7 : fft_fft_SDFChainRadix22__GEN_785; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_787 = 9'hea == fft_fft_SDFChainRadix22__T_215 ? 8'hb8 : fft_fft_SDFChainRadix22__GEN_786; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_788 = 9'heb == fft_fft_SDFChainRadix22__T_215 ? 8'hba : fft_fft_SDFChainRadix22__GEN_787; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_789 = 9'hec == fft_fft_SDFChainRadix22__T_215 ? 8'hbb : fft_fft_SDFChainRadix22__GEN_788; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_790 = 9'hed == fft_fft_SDFChainRadix22__T_215 ? 8'hbc : fft_fft_SDFChainRadix22__GEN_789; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_791 = 9'hee == fft_fft_SDFChainRadix22__T_215 ? 8'hbe : fft_fft_SDFChainRadix22__GEN_790; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_792 = 9'hef == fft_fft_SDFChainRadix22__T_215 ? 8'hbf : fft_fft_SDFChainRadix22__GEN_791; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_793 = 9'hf0 == fft_fft_SDFChainRadix22__T_215 ? 8'hc0 : fft_fft_SDFChainRadix22__GEN_792; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_794 = 9'hf1 == fft_fft_SDFChainRadix22__T_215 ? 8'hc2 : fft_fft_SDFChainRadix22__GEN_793; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_795 = 9'hf2 == fft_fft_SDFChainRadix22__T_215 ? 8'hc3 : fft_fft_SDFChainRadix22__GEN_794; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_796 = 9'hf3 == fft_fft_SDFChainRadix22__T_215 ? 8'hc4 : fft_fft_SDFChainRadix22__GEN_795; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_797 = 9'hf4 == fft_fft_SDFChainRadix22__T_215 ? 8'hc6 : fft_fft_SDFChainRadix22__GEN_796; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_798 = 9'hf5 == fft_fft_SDFChainRadix22__T_215 ? 8'hc7 : fft_fft_SDFChainRadix22__GEN_797; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_799 = 9'hf6 == fft_fft_SDFChainRadix22__T_215 ? 8'hc8 : fft_fft_SDFChainRadix22__GEN_798; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_800 = 9'hf7 == fft_fft_SDFChainRadix22__T_215 ? 8'hca : fft_fft_SDFChainRadix22__GEN_799; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_801 = 9'hf8 == fft_fft_SDFChainRadix22__T_215 ? 8'hcb : fft_fft_SDFChainRadix22__GEN_800; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_802 = 9'hf9 == fft_fft_SDFChainRadix22__T_215 ? 8'hcc : fft_fft_SDFChainRadix22__GEN_801; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_803 = 9'hfa == fft_fft_SDFChainRadix22__T_215 ? 8'hce : fft_fft_SDFChainRadix22__GEN_802; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_804 = 9'hfb == fft_fft_SDFChainRadix22__T_215 ? 8'hcf : fft_fft_SDFChainRadix22__GEN_803; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_805 = 9'hfc == fft_fft_SDFChainRadix22__T_215 ? 8'hd0 : fft_fft_SDFChainRadix22__GEN_804; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_806 = 9'hfd == fft_fft_SDFChainRadix22__T_215 ? 8'hd2 : fft_fft_SDFChainRadix22__GEN_805; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_807 = 9'hfe == fft_fft_SDFChainRadix22__T_215 ? 8'hd3 : fft_fft_SDFChainRadix22__GEN_806; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_808 = 9'hff == fft_fft_SDFChainRadix22__T_215 ? 8'hd4 : fft_fft_SDFChainRadix22__GEN_807; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_809 = 9'h100 == fft_fft_SDFChainRadix22__T_215 ? 8'h0 : fft_fft_SDFChainRadix22__GEN_808; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_810 = 9'h101 == fft_fft_SDFChainRadix22__T_215 ? 8'h1 : fft_fft_SDFChainRadix22__GEN_809; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_811 = 9'h102 == fft_fft_SDFChainRadix22__T_215 ? 8'h2 : fft_fft_SDFChainRadix22__GEN_810; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_812 = 9'h103 == fft_fft_SDFChainRadix22__T_215 ? 8'h3 : fft_fft_SDFChainRadix22__GEN_811; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_813 = 9'h104 == fft_fft_SDFChainRadix22__T_215 ? 8'h4 : fft_fft_SDFChainRadix22__GEN_812; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_814 = 9'h105 == fft_fft_SDFChainRadix22__T_215 ? 8'h5 : fft_fft_SDFChainRadix22__GEN_813; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_815 = 9'h106 == fft_fft_SDFChainRadix22__T_215 ? 8'h6 : fft_fft_SDFChainRadix22__GEN_814; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_816 = 9'h107 == fft_fft_SDFChainRadix22__T_215 ? 8'h7 : fft_fft_SDFChainRadix22__GEN_815; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_817 = 9'h108 == fft_fft_SDFChainRadix22__T_215 ? 8'h8 : fft_fft_SDFChainRadix22__GEN_816; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_818 = 9'h109 == fft_fft_SDFChainRadix22__T_215 ? 8'h9 : fft_fft_SDFChainRadix22__GEN_817; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_819 = 9'h10a == fft_fft_SDFChainRadix22__T_215 ? 8'ha : fft_fft_SDFChainRadix22__GEN_818; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_820 = 9'h10b == fft_fft_SDFChainRadix22__T_215 ? 8'hb : fft_fft_SDFChainRadix22__GEN_819; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_821 = 9'h10c == fft_fft_SDFChainRadix22__T_215 ? 8'hc : fft_fft_SDFChainRadix22__GEN_820; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_822 = 9'h10d == fft_fft_SDFChainRadix22__T_215 ? 8'hd : fft_fft_SDFChainRadix22__GEN_821; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_823 = 9'h10e == fft_fft_SDFChainRadix22__T_215 ? 8'he : fft_fft_SDFChainRadix22__GEN_822; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_824 = 9'h10f == fft_fft_SDFChainRadix22__T_215 ? 8'hf : fft_fft_SDFChainRadix22__GEN_823; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_825 = 9'h110 == fft_fft_SDFChainRadix22__T_215 ? 8'h10 : fft_fft_SDFChainRadix22__GEN_824; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_826 = 9'h111 == fft_fft_SDFChainRadix22__T_215 ? 8'h11 : fft_fft_SDFChainRadix22__GEN_825; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_827 = 9'h112 == fft_fft_SDFChainRadix22__T_215 ? 8'h12 : fft_fft_SDFChainRadix22__GEN_826; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_828 = 9'h113 == fft_fft_SDFChainRadix22__T_215 ? 8'h13 : fft_fft_SDFChainRadix22__GEN_827; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_829 = 9'h114 == fft_fft_SDFChainRadix22__T_215 ? 8'h14 : fft_fft_SDFChainRadix22__GEN_828; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_830 = 9'h115 == fft_fft_SDFChainRadix22__T_215 ? 8'h15 : fft_fft_SDFChainRadix22__GEN_829; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_831 = 9'h116 == fft_fft_SDFChainRadix22__T_215 ? 8'h16 : fft_fft_SDFChainRadix22__GEN_830; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_832 = 9'h117 == fft_fft_SDFChainRadix22__T_215 ? 8'h17 : fft_fft_SDFChainRadix22__GEN_831; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_833 = 9'h118 == fft_fft_SDFChainRadix22__T_215 ? 8'h18 : fft_fft_SDFChainRadix22__GEN_832; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_834 = 9'h119 == fft_fft_SDFChainRadix22__T_215 ? 8'h19 : fft_fft_SDFChainRadix22__GEN_833; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_835 = 9'h11a == fft_fft_SDFChainRadix22__T_215 ? 8'h1a : fft_fft_SDFChainRadix22__GEN_834; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_836 = 9'h11b == fft_fft_SDFChainRadix22__T_215 ? 8'h1b : fft_fft_SDFChainRadix22__GEN_835; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_837 = 9'h11c == fft_fft_SDFChainRadix22__T_215 ? 8'h1c : fft_fft_SDFChainRadix22__GEN_836; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_838 = 9'h11d == fft_fft_SDFChainRadix22__T_215 ? 8'h1d : fft_fft_SDFChainRadix22__GEN_837; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_839 = 9'h11e == fft_fft_SDFChainRadix22__T_215 ? 8'h1e : fft_fft_SDFChainRadix22__GEN_838; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_840 = 9'h11f == fft_fft_SDFChainRadix22__T_215 ? 8'h1f : fft_fft_SDFChainRadix22__GEN_839; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_841 = 9'h120 == fft_fft_SDFChainRadix22__T_215 ? 8'h20 : fft_fft_SDFChainRadix22__GEN_840; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_842 = 9'h121 == fft_fft_SDFChainRadix22__T_215 ? 8'h21 : fft_fft_SDFChainRadix22__GEN_841; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_843 = 9'h122 == fft_fft_SDFChainRadix22__T_215 ? 8'h22 : fft_fft_SDFChainRadix22__GEN_842; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_844 = 9'h123 == fft_fft_SDFChainRadix22__T_215 ? 8'h23 : fft_fft_SDFChainRadix22__GEN_843; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_845 = 9'h124 == fft_fft_SDFChainRadix22__T_215 ? 8'h24 : fft_fft_SDFChainRadix22__GEN_844; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_846 = 9'h125 == fft_fft_SDFChainRadix22__T_215 ? 8'h25 : fft_fft_SDFChainRadix22__GEN_845; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_847 = 9'h126 == fft_fft_SDFChainRadix22__T_215 ? 8'h26 : fft_fft_SDFChainRadix22__GEN_846; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_848 = 9'h127 == fft_fft_SDFChainRadix22__T_215 ? 8'h27 : fft_fft_SDFChainRadix22__GEN_847; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_849 = 9'h128 == fft_fft_SDFChainRadix22__T_215 ? 8'h28 : fft_fft_SDFChainRadix22__GEN_848; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_850 = 9'h129 == fft_fft_SDFChainRadix22__T_215 ? 8'h29 : fft_fft_SDFChainRadix22__GEN_849; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_851 = 9'h12a == fft_fft_SDFChainRadix22__T_215 ? 8'h2a : fft_fft_SDFChainRadix22__GEN_850; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_852 = 9'h12b == fft_fft_SDFChainRadix22__T_215 ? 8'h2b : fft_fft_SDFChainRadix22__GEN_851; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_853 = 9'h12c == fft_fft_SDFChainRadix22__T_215 ? 8'h2c : fft_fft_SDFChainRadix22__GEN_852; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_854 = 9'h12d == fft_fft_SDFChainRadix22__T_215 ? 8'h2d : fft_fft_SDFChainRadix22__GEN_853; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_855 = 9'h12e == fft_fft_SDFChainRadix22__T_215 ? 8'h2e : fft_fft_SDFChainRadix22__GEN_854; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_856 = 9'h12f == fft_fft_SDFChainRadix22__T_215 ? 8'h2f : fft_fft_SDFChainRadix22__GEN_855; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_857 = 9'h130 == fft_fft_SDFChainRadix22__T_215 ? 8'h30 : fft_fft_SDFChainRadix22__GEN_856; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_858 = 9'h131 == fft_fft_SDFChainRadix22__T_215 ? 8'h31 : fft_fft_SDFChainRadix22__GEN_857; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_859 = 9'h132 == fft_fft_SDFChainRadix22__T_215 ? 8'h32 : fft_fft_SDFChainRadix22__GEN_858; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_860 = 9'h133 == fft_fft_SDFChainRadix22__T_215 ? 8'h33 : fft_fft_SDFChainRadix22__GEN_859; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_861 = 9'h134 == fft_fft_SDFChainRadix22__T_215 ? 8'h34 : fft_fft_SDFChainRadix22__GEN_860; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_862 = 9'h135 == fft_fft_SDFChainRadix22__T_215 ? 8'h35 : fft_fft_SDFChainRadix22__GEN_861; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_863 = 9'h136 == fft_fft_SDFChainRadix22__T_215 ? 8'h36 : fft_fft_SDFChainRadix22__GEN_862; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_864 = 9'h137 == fft_fft_SDFChainRadix22__T_215 ? 8'h37 : fft_fft_SDFChainRadix22__GEN_863; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_865 = 9'h138 == fft_fft_SDFChainRadix22__T_215 ? 8'h38 : fft_fft_SDFChainRadix22__GEN_864; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_866 = 9'h139 == fft_fft_SDFChainRadix22__T_215 ? 8'h39 : fft_fft_SDFChainRadix22__GEN_865; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_867 = 9'h13a == fft_fft_SDFChainRadix22__T_215 ? 8'h3a : fft_fft_SDFChainRadix22__GEN_866; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_868 = 9'h13b == fft_fft_SDFChainRadix22__T_215 ? 8'h3b : fft_fft_SDFChainRadix22__GEN_867; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_869 = 9'h13c == fft_fft_SDFChainRadix22__T_215 ? 8'h3c : fft_fft_SDFChainRadix22__GEN_868; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_870 = 9'h13d == fft_fft_SDFChainRadix22__T_215 ? 8'h3d : fft_fft_SDFChainRadix22__GEN_869; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_871 = 9'h13e == fft_fft_SDFChainRadix22__T_215 ? 8'h3e : fft_fft_SDFChainRadix22__GEN_870; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_872 = 9'h13f == fft_fft_SDFChainRadix22__T_215 ? 8'h3f : fft_fft_SDFChainRadix22__GEN_871; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_873 = 9'h140 == fft_fft_SDFChainRadix22__T_215 ? 8'h40 : fft_fft_SDFChainRadix22__GEN_872; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_874 = 9'h141 == fft_fft_SDFChainRadix22__T_215 ? 8'h41 : fft_fft_SDFChainRadix22__GEN_873; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_875 = 9'h142 == fft_fft_SDFChainRadix22__T_215 ? 8'h42 : fft_fft_SDFChainRadix22__GEN_874; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_876 = 9'h143 == fft_fft_SDFChainRadix22__T_215 ? 8'h43 : fft_fft_SDFChainRadix22__GEN_875; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_877 = 9'h144 == fft_fft_SDFChainRadix22__T_215 ? 8'h44 : fft_fft_SDFChainRadix22__GEN_876; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_878 = 9'h145 == fft_fft_SDFChainRadix22__T_215 ? 8'h45 : fft_fft_SDFChainRadix22__GEN_877; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_879 = 9'h146 == fft_fft_SDFChainRadix22__T_215 ? 8'h46 : fft_fft_SDFChainRadix22__GEN_878; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_880 = 9'h147 == fft_fft_SDFChainRadix22__T_215 ? 8'h47 : fft_fft_SDFChainRadix22__GEN_879; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_881 = 9'h148 == fft_fft_SDFChainRadix22__T_215 ? 8'h48 : fft_fft_SDFChainRadix22__GEN_880; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_882 = 9'h149 == fft_fft_SDFChainRadix22__T_215 ? 8'h49 : fft_fft_SDFChainRadix22__GEN_881; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_883 = 9'h14a == fft_fft_SDFChainRadix22__T_215 ? 8'h4a : fft_fft_SDFChainRadix22__GEN_882; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_884 = 9'h14b == fft_fft_SDFChainRadix22__T_215 ? 8'h4b : fft_fft_SDFChainRadix22__GEN_883; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_885 = 9'h14c == fft_fft_SDFChainRadix22__T_215 ? 8'h4c : fft_fft_SDFChainRadix22__GEN_884; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_886 = 9'h14d == fft_fft_SDFChainRadix22__T_215 ? 8'h4d : fft_fft_SDFChainRadix22__GEN_885; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_887 = 9'h14e == fft_fft_SDFChainRadix22__T_215 ? 8'h4e : fft_fft_SDFChainRadix22__GEN_886; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_888 = 9'h14f == fft_fft_SDFChainRadix22__T_215 ? 8'h4f : fft_fft_SDFChainRadix22__GEN_887; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_889 = 9'h150 == fft_fft_SDFChainRadix22__T_215 ? 8'h50 : fft_fft_SDFChainRadix22__GEN_888; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_890 = 9'h151 == fft_fft_SDFChainRadix22__T_215 ? 8'h51 : fft_fft_SDFChainRadix22__GEN_889; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_891 = 9'h152 == fft_fft_SDFChainRadix22__T_215 ? 8'h52 : fft_fft_SDFChainRadix22__GEN_890; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_892 = 9'h153 == fft_fft_SDFChainRadix22__T_215 ? 8'h53 : fft_fft_SDFChainRadix22__GEN_891; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_893 = 9'h154 == fft_fft_SDFChainRadix22__T_215 ? 8'h54 : fft_fft_SDFChainRadix22__GEN_892; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_894 = 9'h155 == fft_fft_SDFChainRadix22__T_215 ? 8'h55 : fft_fft_SDFChainRadix22__GEN_893; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_895 = 9'h156 == fft_fft_SDFChainRadix22__T_215 ? 8'h56 : fft_fft_SDFChainRadix22__GEN_894; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_896 = 9'h157 == fft_fft_SDFChainRadix22__T_215 ? 8'h57 : fft_fft_SDFChainRadix22__GEN_895; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_897 = 9'h158 == fft_fft_SDFChainRadix22__T_215 ? 8'h58 : fft_fft_SDFChainRadix22__GEN_896; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_898 = 9'h159 == fft_fft_SDFChainRadix22__T_215 ? 8'h59 : fft_fft_SDFChainRadix22__GEN_897; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_899 = 9'h15a == fft_fft_SDFChainRadix22__T_215 ? 8'h5a : fft_fft_SDFChainRadix22__GEN_898; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_900 = 9'h15b == fft_fft_SDFChainRadix22__T_215 ? 8'h5b : fft_fft_SDFChainRadix22__GEN_899; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_901 = 9'h15c == fft_fft_SDFChainRadix22__T_215 ? 8'h5c : fft_fft_SDFChainRadix22__GEN_900; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_902 = 9'h15d == fft_fft_SDFChainRadix22__T_215 ? 8'h5d : fft_fft_SDFChainRadix22__GEN_901; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_903 = 9'h15e == fft_fft_SDFChainRadix22__T_215 ? 8'h5e : fft_fft_SDFChainRadix22__GEN_902; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_904 = 9'h15f == fft_fft_SDFChainRadix22__T_215 ? 8'h5f : fft_fft_SDFChainRadix22__GEN_903; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_905 = 9'h160 == fft_fft_SDFChainRadix22__T_215 ? 8'h60 : fft_fft_SDFChainRadix22__GEN_904; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_906 = 9'h161 == fft_fft_SDFChainRadix22__T_215 ? 8'h61 : fft_fft_SDFChainRadix22__GEN_905; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_907 = 9'h162 == fft_fft_SDFChainRadix22__T_215 ? 8'h62 : fft_fft_SDFChainRadix22__GEN_906; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_908 = 9'h163 == fft_fft_SDFChainRadix22__T_215 ? 8'h63 : fft_fft_SDFChainRadix22__GEN_907; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_909 = 9'h164 == fft_fft_SDFChainRadix22__T_215 ? 8'h64 : fft_fft_SDFChainRadix22__GEN_908; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_910 = 9'h165 == fft_fft_SDFChainRadix22__T_215 ? 8'h65 : fft_fft_SDFChainRadix22__GEN_909; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_911 = 9'h166 == fft_fft_SDFChainRadix22__T_215 ? 8'h66 : fft_fft_SDFChainRadix22__GEN_910; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_912 = 9'h167 == fft_fft_SDFChainRadix22__T_215 ? 8'h67 : fft_fft_SDFChainRadix22__GEN_911; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_913 = 9'h168 == fft_fft_SDFChainRadix22__T_215 ? 8'h68 : fft_fft_SDFChainRadix22__GEN_912; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_914 = 9'h169 == fft_fft_SDFChainRadix22__T_215 ? 8'h69 : fft_fft_SDFChainRadix22__GEN_913; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_915 = 9'h16a == fft_fft_SDFChainRadix22__T_215 ? 8'h6a : fft_fft_SDFChainRadix22__GEN_914; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_916 = 9'h16b == fft_fft_SDFChainRadix22__T_215 ? 8'h6b : fft_fft_SDFChainRadix22__GEN_915; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_917 = 9'h16c == fft_fft_SDFChainRadix22__T_215 ? 8'h6c : fft_fft_SDFChainRadix22__GEN_916; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_918 = 9'h16d == fft_fft_SDFChainRadix22__T_215 ? 8'h6d : fft_fft_SDFChainRadix22__GEN_917; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_919 = 9'h16e == fft_fft_SDFChainRadix22__T_215 ? 8'h6e : fft_fft_SDFChainRadix22__GEN_918; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_920 = 9'h16f == fft_fft_SDFChainRadix22__T_215 ? 8'h6f : fft_fft_SDFChainRadix22__GEN_919; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_921 = 9'h170 == fft_fft_SDFChainRadix22__T_215 ? 8'h70 : fft_fft_SDFChainRadix22__GEN_920; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_922 = 9'h171 == fft_fft_SDFChainRadix22__T_215 ? 8'h71 : fft_fft_SDFChainRadix22__GEN_921; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_923 = 9'h172 == fft_fft_SDFChainRadix22__T_215 ? 8'h72 : fft_fft_SDFChainRadix22__GEN_922; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_924 = 9'h173 == fft_fft_SDFChainRadix22__T_215 ? 8'h73 : fft_fft_SDFChainRadix22__GEN_923; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_925 = 9'h174 == fft_fft_SDFChainRadix22__T_215 ? 8'h74 : fft_fft_SDFChainRadix22__GEN_924; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_926 = 9'h175 == fft_fft_SDFChainRadix22__T_215 ? 8'h75 : fft_fft_SDFChainRadix22__GEN_925; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_927 = 9'h176 == fft_fft_SDFChainRadix22__T_215 ? 8'h76 : fft_fft_SDFChainRadix22__GEN_926; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_928 = 9'h177 == fft_fft_SDFChainRadix22__T_215 ? 8'h77 : fft_fft_SDFChainRadix22__GEN_927; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_929 = 9'h178 == fft_fft_SDFChainRadix22__T_215 ? 8'h78 : fft_fft_SDFChainRadix22__GEN_928; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_930 = 9'h179 == fft_fft_SDFChainRadix22__T_215 ? 8'h79 : fft_fft_SDFChainRadix22__GEN_929; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_931 = 9'h17a == fft_fft_SDFChainRadix22__T_215 ? 8'h7a : fft_fft_SDFChainRadix22__GEN_930; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_932 = 9'h17b == fft_fft_SDFChainRadix22__T_215 ? 8'h7b : fft_fft_SDFChainRadix22__GEN_931; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_933 = 9'h17c == fft_fft_SDFChainRadix22__T_215 ? 8'h7c : fft_fft_SDFChainRadix22__GEN_932; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_934 = 9'h17d == fft_fft_SDFChainRadix22__T_215 ? 8'h7d : fft_fft_SDFChainRadix22__GEN_933; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_935 = 9'h17e == fft_fft_SDFChainRadix22__T_215 ? 8'h7e : fft_fft_SDFChainRadix22__GEN_934; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_936 = 9'h17f == fft_fft_SDFChainRadix22__T_215 ? 8'h7f : fft_fft_SDFChainRadix22__GEN_935; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_937 = 9'h180 == fft_fft_SDFChainRadix22__T_215 ? 8'h0 : fft_fft_SDFChainRadix22__GEN_936; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_938 = 9'h181 == fft_fft_SDFChainRadix22__T_215 ? 8'h3 : fft_fft_SDFChainRadix22__GEN_937; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_939 = 9'h182 == fft_fft_SDFChainRadix22__T_215 ? 8'h6 : fft_fft_SDFChainRadix22__GEN_938; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_940 = 9'h183 == fft_fft_SDFChainRadix22__T_215 ? 8'h9 : fft_fft_SDFChainRadix22__GEN_939; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_941 = 9'h184 == fft_fft_SDFChainRadix22__T_215 ? 8'hc : fft_fft_SDFChainRadix22__GEN_940; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_942 = 9'h185 == fft_fft_SDFChainRadix22__T_215 ? 8'hf : fft_fft_SDFChainRadix22__GEN_941; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_943 = 9'h186 == fft_fft_SDFChainRadix22__T_215 ? 8'h12 : fft_fft_SDFChainRadix22__GEN_942; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_944 = 9'h187 == fft_fft_SDFChainRadix22__T_215 ? 8'h15 : fft_fft_SDFChainRadix22__GEN_943; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_945 = 9'h188 == fft_fft_SDFChainRadix22__T_215 ? 8'h18 : fft_fft_SDFChainRadix22__GEN_944; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_946 = 9'h189 == fft_fft_SDFChainRadix22__T_215 ? 8'h1b : fft_fft_SDFChainRadix22__GEN_945; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_947 = 9'h18a == fft_fft_SDFChainRadix22__T_215 ? 8'h1e : fft_fft_SDFChainRadix22__GEN_946; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_948 = 9'h18b == fft_fft_SDFChainRadix22__T_215 ? 8'h21 : fft_fft_SDFChainRadix22__GEN_947; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_949 = 9'h18c == fft_fft_SDFChainRadix22__T_215 ? 8'h24 : fft_fft_SDFChainRadix22__GEN_948; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_950 = 9'h18d == fft_fft_SDFChainRadix22__T_215 ? 8'h27 : fft_fft_SDFChainRadix22__GEN_949; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_951 = 9'h18e == fft_fft_SDFChainRadix22__T_215 ? 8'h2a : fft_fft_SDFChainRadix22__GEN_950; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_952 = 9'h18f == fft_fft_SDFChainRadix22__T_215 ? 8'h2d : fft_fft_SDFChainRadix22__GEN_951; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_953 = 9'h190 == fft_fft_SDFChainRadix22__T_215 ? 8'h30 : fft_fft_SDFChainRadix22__GEN_952; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_954 = 9'h191 == fft_fft_SDFChainRadix22__T_215 ? 8'h33 : fft_fft_SDFChainRadix22__GEN_953; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_955 = 9'h192 == fft_fft_SDFChainRadix22__T_215 ? 8'h36 : fft_fft_SDFChainRadix22__GEN_954; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_956 = 9'h193 == fft_fft_SDFChainRadix22__T_215 ? 8'h39 : fft_fft_SDFChainRadix22__GEN_955; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_957 = 9'h194 == fft_fft_SDFChainRadix22__T_215 ? 8'h3c : fft_fft_SDFChainRadix22__GEN_956; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_958 = 9'h195 == fft_fft_SDFChainRadix22__T_215 ? 8'h3f : fft_fft_SDFChainRadix22__GEN_957; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_959 = 9'h196 == fft_fft_SDFChainRadix22__T_215 ? 8'h42 : fft_fft_SDFChainRadix22__GEN_958; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_960 = 9'h197 == fft_fft_SDFChainRadix22__T_215 ? 8'h45 : fft_fft_SDFChainRadix22__GEN_959; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_961 = 9'h198 == fft_fft_SDFChainRadix22__T_215 ? 8'h48 : fft_fft_SDFChainRadix22__GEN_960; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_962 = 9'h199 == fft_fft_SDFChainRadix22__T_215 ? 8'h4b : fft_fft_SDFChainRadix22__GEN_961; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_963 = 9'h19a == fft_fft_SDFChainRadix22__T_215 ? 8'h4e : fft_fft_SDFChainRadix22__GEN_962; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_964 = 9'h19b == fft_fft_SDFChainRadix22__T_215 ? 8'h51 : fft_fft_SDFChainRadix22__GEN_963; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_965 = 9'h19c == fft_fft_SDFChainRadix22__T_215 ? 8'h54 : fft_fft_SDFChainRadix22__GEN_964; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_966 = 9'h19d == fft_fft_SDFChainRadix22__T_215 ? 8'h57 : fft_fft_SDFChainRadix22__GEN_965; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_967 = 9'h19e == fft_fft_SDFChainRadix22__T_215 ? 8'h5a : fft_fft_SDFChainRadix22__GEN_966; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_968 = 9'h19f == fft_fft_SDFChainRadix22__T_215 ? 8'h5d : fft_fft_SDFChainRadix22__GEN_967; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_969 = 9'h1a0 == fft_fft_SDFChainRadix22__T_215 ? 8'h60 : fft_fft_SDFChainRadix22__GEN_968; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_970 = 9'h1a1 == fft_fft_SDFChainRadix22__T_215 ? 8'h63 : fft_fft_SDFChainRadix22__GEN_969; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_971 = 9'h1a2 == fft_fft_SDFChainRadix22__T_215 ? 8'h66 : fft_fft_SDFChainRadix22__GEN_970; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_972 = 9'h1a3 == fft_fft_SDFChainRadix22__T_215 ? 8'h69 : fft_fft_SDFChainRadix22__GEN_971; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_973 = 9'h1a4 == fft_fft_SDFChainRadix22__T_215 ? 8'h6c : fft_fft_SDFChainRadix22__GEN_972; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_974 = 9'h1a5 == fft_fft_SDFChainRadix22__T_215 ? 8'h6f : fft_fft_SDFChainRadix22__GEN_973; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_975 = 9'h1a6 == fft_fft_SDFChainRadix22__T_215 ? 8'h72 : fft_fft_SDFChainRadix22__GEN_974; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_976 = 9'h1a7 == fft_fft_SDFChainRadix22__T_215 ? 8'h75 : fft_fft_SDFChainRadix22__GEN_975; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_977 = 9'h1a8 == fft_fft_SDFChainRadix22__T_215 ? 8'h78 : fft_fft_SDFChainRadix22__GEN_976; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_978 = 9'h1a9 == fft_fft_SDFChainRadix22__T_215 ? 8'h7b : fft_fft_SDFChainRadix22__GEN_977; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_979 = 9'h1aa == fft_fft_SDFChainRadix22__T_215 ? 8'h7e : fft_fft_SDFChainRadix22__GEN_978; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_980 = 9'h1ab == fft_fft_SDFChainRadix22__T_215 ? 8'h81 : fft_fft_SDFChainRadix22__GEN_979; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_981 = 9'h1ac == fft_fft_SDFChainRadix22__T_215 ? 8'h83 : fft_fft_SDFChainRadix22__GEN_980; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_982 = 9'h1ad == fft_fft_SDFChainRadix22__T_215 ? 8'h85 : fft_fft_SDFChainRadix22__GEN_981; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_983 = 9'h1ae == fft_fft_SDFChainRadix22__T_215 ? 8'h87 : fft_fft_SDFChainRadix22__GEN_982; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_984 = 9'h1af == fft_fft_SDFChainRadix22__T_215 ? 8'h89 : fft_fft_SDFChainRadix22__GEN_983; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_985 = 9'h1b0 == fft_fft_SDFChainRadix22__T_215 ? 8'h8b : fft_fft_SDFChainRadix22__GEN_984; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_986 = 9'h1b1 == fft_fft_SDFChainRadix22__T_215 ? 8'h8d : fft_fft_SDFChainRadix22__GEN_985; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_987 = 9'h1b2 == fft_fft_SDFChainRadix22__T_215 ? 8'h8f : fft_fft_SDFChainRadix22__GEN_986; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_988 = 9'h1b3 == fft_fft_SDFChainRadix22__T_215 ? 8'h91 : fft_fft_SDFChainRadix22__GEN_987; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_989 = 9'h1b4 == fft_fft_SDFChainRadix22__T_215 ? 8'h93 : fft_fft_SDFChainRadix22__GEN_988; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_990 = 9'h1b5 == fft_fft_SDFChainRadix22__T_215 ? 8'h95 : fft_fft_SDFChainRadix22__GEN_989; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_991 = 9'h1b6 == fft_fft_SDFChainRadix22__T_215 ? 8'h97 : fft_fft_SDFChainRadix22__GEN_990; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_992 = 9'h1b7 == fft_fft_SDFChainRadix22__T_215 ? 8'h99 : fft_fft_SDFChainRadix22__GEN_991; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_993 = 9'h1b8 == fft_fft_SDFChainRadix22__T_215 ? 8'h9b : fft_fft_SDFChainRadix22__GEN_992; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_994 = 9'h1b9 == fft_fft_SDFChainRadix22__T_215 ? 8'h9d : fft_fft_SDFChainRadix22__GEN_993; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_995 = 9'h1ba == fft_fft_SDFChainRadix22__T_215 ? 8'h9f : fft_fft_SDFChainRadix22__GEN_994; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_996 = 9'h1bb == fft_fft_SDFChainRadix22__T_215 ? 8'ha1 : fft_fft_SDFChainRadix22__GEN_995; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_997 = 9'h1bc == fft_fft_SDFChainRadix22__T_215 ? 8'ha3 : fft_fft_SDFChainRadix22__GEN_996; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_998 = 9'h1bd == fft_fft_SDFChainRadix22__T_215 ? 8'ha5 : fft_fft_SDFChainRadix22__GEN_997; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_999 = 9'h1be == fft_fft_SDFChainRadix22__T_215 ? 8'ha7 : fft_fft_SDFChainRadix22__GEN_998; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1000 = 9'h1bf == fft_fft_SDFChainRadix22__T_215 ? 8'ha9 : fft_fft_SDFChainRadix22__GEN_999; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1001 = 9'h1c0 == fft_fft_SDFChainRadix22__T_215 ? 8'hab : fft_fft_SDFChainRadix22__GEN_1000; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1002 = 9'h1c1 == fft_fft_SDFChainRadix22__T_215 ? 8'had : fft_fft_SDFChainRadix22__GEN_1001; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1003 = 9'h1c2 == fft_fft_SDFChainRadix22__T_215 ? 8'haf : fft_fft_SDFChainRadix22__GEN_1002; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1004 = 9'h1c3 == fft_fft_SDFChainRadix22__T_215 ? 8'hb1 : fft_fft_SDFChainRadix22__GEN_1003; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1005 = 9'h1c4 == fft_fft_SDFChainRadix22__T_215 ? 8'hb3 : fft_fft_SDFChainRadix22__GEN_1004; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1006 = 9'h1c5 == fft_fft_SDFChainRadix22__T_215 ? 8'hb5 : fft_fft_SDFChainRadix22__GEN_1005; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1007 = 9'h1c6 == fft_fft_SDFChainRadix22__T_215 ? 8'hb7 : fft_fft_SDFChainRadix22__GEN_1006; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1008 = 9'h1c7 == fft_fft_SDFChainRadix22__T_215 ? 8'hb9 : fft_fft_SDFChainRadix22__GEN_1007; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1009 = 9'h1c8 == fft_fft_SDFChainRadix22__T_215 ? 8'hbb : fft_fft_SDFChainRadix22__GEN_1008; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1010 = 9'h1c9 == fft_fft_SDFChainRadix22__T_215 ? 8'hbd : fft_fft_SDFChainRadix22__GEN_1009; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1011 = 9'h1ca == fft_fft_SDFChainRadix22__T_215 ? 8'hbf : fft_fft_SDFChainRadix22__GEN_1010; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1012 = 9'h1cb == fft_fft_SDFChainRadix22__T_215 ? 8'hc1 : fft_fft_SDFChainRadix22__GEN_1011; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1013 = 9'h1cc == fft_fft_SDFChainRadix22__T_215 ? 8'hc3 : fft_fft_SDFChainRadix22__GEN_1012; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1014 = 9'h1cd == fft_fft_SDFChainRadix22__T_215 ? 8'hc5 : fft_fft_SDFChainRadix22__GEN_1013; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1015 = 9'h1ce == fft_fft_SDFChainRadix22__T_215 ? 8'hc7 : fft_fft_SDFChainRadix22__GEN_1014; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1016 = 9'h1cf == fft_fft_SDFChainRadix22__T_215 ? 8'hc9 : fft_fft_SDFChainRadix22__GEN_1015; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1017 = 9'h1d0 == fft_fft_SDFChainRadix22__T_215 ? 8'hcb : fft_fft_SDFChainRadix22__GEN_1016; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1018 = 9'h1d1 == fft_fft_SDFChainRadix22__T_215 ? 8'hcd : fft_fft_SDFChainRadix22__GEN_1017; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1019 = 9'h1d2 == fft_fft_SDFChainRadix22__T_215 ? 8'hcf : fft_fft_SDFChainRadix22__GEN_1018; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1020 = 9'h1d3 == fft_fft_SDFChainRadix22__T_215 ? 8'hd1 : fft_fft_SDFChainRadix22__GEN_1019; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1021 = 9'h1d4 == fft_fft_SDFChainRadix22__T_215 ? 8'hd3 : fft_fft_SDFChainRadix22__GEN_1020; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1022 = 9'h1d5 == fft_fft_SDFChainRadix22__T_215 ? 8'hd5 : fft_fft_SDFChainRadix22__GEN_1021; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1023 = 9'h1d6 == fft_fft_SDFChainRadix22__T_215 ? 8'hd6 : fft_fft_SDFChainRadix22__GEN_1022; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1024 = 9'h1d7 == fft_fft_SDFChainRadix22__T_215 ? 8'hd7 : fft_fft_SDFChainRadix22__GEN_1023; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1025 = 9'h1d8 == fft_fft_SDFChainRadix22__T_215 ? 8'hd8 : fft_fft_SDFChainRadix22__GEN_1024; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1026 = 9'h1d9 == fft_fft_SDFChainRadix22__T_215 ? 8'hd9 : fft_fft_SDFChainRadix22__GEN_1025; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1027 = 9'h1da == fft_fft_SDFChainRadix22__T_215 ? 8'hda : fft_fft_SDFChainRadix22__GEN_1026; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1028 = 9'h1db == fft_fft_SDFChainRadix22__T_215 ? 8'hdb : fft_fft_SDFChainRadix22__GEN_1027; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1029 = 9'h1dc == fft_fft_SDFChainRadix22__T_215 ? 8'hdc : fft_fft_SDFChainRadix22__GEN_1028; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1030 = 9'h1dd == fft_fft_SDFChainRadix22__T_215 ? 8'hdd : fft_fft_SDFChainRadix22__GEN_1029; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1031 = 9'h1de == fft_fft_SDFChainRadix22__T_215 ? 8'hde : fft_fft_SDFChainRadix22__GEN_1030; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1032 = 9'h1df == fft_fft_SDFChainRadix22__T_215 ? 8'hdf : fft_fft_SDFChainRadix22__GEN_1031; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1033 = 9'h1e0 == fft_fft_SDFChainRadix22__T_215 ? 8'he0 : fft_fft_SDFChainRadix22__GEN_1032; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1034 = 9'h1e1 == fft_fft_SDFChainRadix22__T_215 ? 8'he1 : fft_fft_SDFChainRadix22__GEN_1033; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1035 = 9'h1e2 == fft_fft_SDFChainRadix22__T_215 ? 8'he2 : fft_fft_SDFChainRadix22__GEN_1034; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1036 = 9'h1e3 == fft_fft_SDFChainRadix22__T_215 ? 8'he3 : fft_fft_SDFChainRadix22__GEN_1035; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1037 = 9'h1e4 == fft_fft_SDFChainRadix22__T_215 ? 8'he4 : fft_fft_SDFChainRadix22__GEN_1036; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1038 = 9'h1e5 == fft_fft_SDFChainRadix22__T_215 ? 8'he5 : fft_fft_SDFChainRadix22__GEN_1037; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1039 = 9'h1e6 == fft_fft_SDFChainRadix22__T_215 ? 8'he6 : fft_fft_SDFChainRadix22__GEN_1038; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1040 = 9'h1e7 == fft_fft_SDFChainRadix22__T_215 ? 8'he7 : fft_fft_SDFChainRadix22__GEN_1039; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1041 = 9'h1e8 == fft_fft_SDFChainRadix22__T_215 ? 8'he8 : fft_fft_SDFChainRadix22__GEN_1040; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1042 = 9'h1e9 == fft_fft_SDFChainRadix22__T_215 ? 8'he9 : fft_fft_SDFChainRadix22__GEN_1041; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1043 = 9'h1ea == fft_fft_SDFChainRadix22__T_215 ? 8'hea : fft_fft_SDFChainRadix22__GEN_1042; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1044 = 9'h1eb == fft_fft_SDFChainRadix22__T_215 ? 8'heb : fft_fft_SDFChainRadix22__GEN_1043; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1045 = 9'h1ec == fft_fft_SDFChainRadix22__T_215 ? 8'hec : fft_fft_SDFChainRadix22__GEN_1044; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1046 = 9'h1ed == fft_fft_SDFChainRadix22__T_215 ? 8'hed : fft_fft_SDFChainRadix22__GEN_1045; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1047 = 9'h1ee == fft_fft_SDFChainRadix22__T_215 ? 8'hee : fft_fft_SDFChainRadix22__GEN_1046; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1048 = 9'h1ef == fft_fft_SDFChainRadix22__T_215 ? 8'hef : fft_fft_SDFChainRadix22__GEN_1047; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1049 = 9'h1f0 == fft_fft_SDFChainRadix22__T_215 ? 8'hf0 : fft_fft_SDFChainRadix22__GEN_1048; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1050 = 9'h1f1 == fft_fft_SDFChainRadix22__T_215 ? 8'hf1 : fft_fft_SDFChainRadix22__GEN_1049; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1051 = 9'h1f2 == fft_fft_SDFChainRadix22__T_215 ? 8'hf2 : fft_fft_SDFChainRadix22__GEN_1050; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1052 = 9'h1f3 == fft_fft_SDFChainRadix22__T_215 ? 8'hf3 : fft_fft_SDFChainRadix22__GEN_1051; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1053 = 9'h1f4 == fft_fft_SDFChainRadix22__T_215 ? 8'hf4 : fft_fft_SDFChainRadix22__GEN_1052; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1054 = 9'h1f5 == fft_fft_SDFChainRadix22__T_215 ? 8'hf5 : fft_fft_SDFChainRadix22__GEN_1053; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1055 = 9'h1f6 == fft_fft_SDFChainRadix22__T_215 ? 8'hf6 : fft_fft_SDFChainRadix22__GEN_1054; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1056 = 9'h1f7 == fft_fft_SDFChainRadix22__T_215 ? 8'hf7 : fft_fft_SDFChainRadix22__GEN_1055; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1057 = 9'h1f8 == fft_fft_SDFChainRadix22__T_215 ? 8'hf8 : fft_fft_SDFChainRadix22__GEN_1056; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1058 = 9'h1f9 == fft_fft_SDFChainRadix22__T_215 ? 8'hf9 : fft_fft_SDFChainRadix22__GEN_1057; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1059 = 9'h1fa == fft_fft_SDFChainRadix22__T_215 ? 8'hfa : fft_fft_SDFChainRadix22__GEN_1058; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1060 = 9'h1fb == fft_fft_SDFChainRadix22__T_215 ? 8'hfb : fft_fft_SDFChainRadix22__GEN_1059; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1061 = 9'h1fc == fft_fft_SDFChainRadix22__T_215 ? 8'hfc : fft_fft_SDFChainRadix22__GEN_1060; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1062 = 9'h1fd == fft_fft_SDFChainRadix22__T_215 ? 8'hfd : fft_fft_SDFChainRadix22__GEN_1061; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1063 = 9'h1fe == fft_fft_SDFChainRadix22__T_215 ? 8'hfe : fft_fft_SDFChainRadix22__GEN_1062; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1064 = 9'h1ff == fft_fft_SDFChainRadix22__T_215 ? 8'hff : fft_fft_SDFChainRadix22__GEN_1063; // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1067 = 8'h1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3fff) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1068 = 8'h1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shc9) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1069 = 8'h2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ffb) : $signed(fft_fft_SDFChainRadix22__GEN_1067); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1070 = 8'h2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh192) : $signed(fft_fft_SDFChainRadix22__GEN_1068); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1071 = 8'h3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ff5) : $signed(fft_fft_SDFChainRadix22__GEN_1069); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1072 = 8'h3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh25b) : $signed(fft_fft_SDFChainRadix22__GEN_1070); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1073 = 8'h4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3fec) : $signed(fft_fft_SDFChainRadix22__GEN_1071); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1074 = 8'h4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh324) : $signed(fft_fft_SDFChainRadix22__GEN_1072); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1075 = 8'h5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3fe1) : $signed(fft_fft_SDFChainRadix22__GEN_1073); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1076 = 8'h5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ed) : $signed(fft_fft_SDFChainRadix22__GEN_1074); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1077 = 8'h6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3fd4) : $signed(fft_fft_SDFChainRadix22__GEN_1075); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1078 = 8'h6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh4b5) : $signed(fft_fft_SDFChainRadix22__GEN_1076); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1079 = 8'h7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3fc4) : $signed(fft_fft_SDFChainRadix22__GEN_1077); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1080 = 8'h7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh57e) : $signed(fft_fft_SDFChainRadix22__GEN_1078); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1081 = 8'h8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_1079); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1082 = 8'h8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_1080); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1083 = 8'h9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f9c) : $signed(fft_fft_SDFChainRadix22__GEN_1081); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1084 = 8'h9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh70e) : $signed(fft_fft_SDFChainRadix22__GEN_1082); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1085 = 8'ha == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f85) : $signed(fft_fft_SDFChainRadix22__GEN_1083); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1086 = 8'ha == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh7d6) : $signed(fft_fft_SDFChainRadix22__GEN_1084); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1087 = 8'hb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f6b) : $signed(fft_fft_SDFChainRadix22__GEN_1085); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1088 = 8'hb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh89d) : $signed(fft_fft_SDFChainRadix22__GEN_1086); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1089 = 8'hc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_1087); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1090 = 8'hc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_1088); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1091 = 8'hd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f30) : $signed(fft_fft_SDFChainRadix22__GEN_1089); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1092 = 8'hd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sha2b) : $signed(fft_fft_SDFChainRadix22__GEN_1090); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1093 = 8'he == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f0f) : $signed(fft_fft_SDFChainRadix22__GEN_1091); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1094 = 8'he == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shaf1) : $signed(fft_fft_SDFChainRadix22__GEN_1092); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1095 = 8'hf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3eeb) : $signed(fft_fft_SDFChainRadix22__GEN_1093); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1096 = 8'hf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shbb7) : $signed(fft_fft_SDFChainRadix22__GEN_1094); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1097 = 8'h10 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_1095); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1098 = 8'h10 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_1096); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1099 = 8'h11 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3e9d) : $signed(fft_fft_SDFChainRadix22__GEN_1097); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1100 = 8'h11 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shd41) : $signed(fft_fft_SDFChainRadix22__GEN_1098); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1101 = 8'h12 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3e72) : $signed(fft_fft_SDFChainRadix22__GEN_1099); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1102 = 8'h12 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'she06) : $signed(fft_fft_SDFChainRadix22__GEN_1100); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1103 = 8'h13 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3e45) : $signed(fft_fft_SDFChainRadix22__GEN_1101); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1104 = 8'h13 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sheca) : $signed(fft_fft_SDFChainRadix22__GEN_1102); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1105 = 8'h14 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_1103); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1106 = 8'h14 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_1104); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1107 = 8'h15 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3de3) : $signed(fft_fft_SDFChainRadix22__GEN_1105); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1108 = 8'h15 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1050) : $signed(fft_fft_SDFChainRadix22__GEN_1106); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1109 = 8'h16 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3daf) : $signed(fft_fft_SDFChainRadix22__GEN_1107); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1110 = 8'h16 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1112) : $signed(fft_fft_SDFChainRadix22__GEN_1108); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1111 = 8'h17 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3d78) : $signed(fft_fft_SDFChainRadix22__GEN_1109); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1112 = 8'h17 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh11d3) : $signed(fft_fft_SDFChainRadix22__GEN_1110); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1113 = 8'h18 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_1111); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1114 = 8'h18 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_1112); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1115 = 8'h19 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3d03) : $signed(fft_fft_SDFChainRadix22__GEN_1113); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1116 = 8'h19 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1354) : $signed(fft_fft_SDFChainRadix22__GEN_1114); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1117 = 8'h1a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3cc5) : $signed(fft_fft_SDFChainRadix22__GEN_1115); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1118 = 8'h1a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1413) : $signed(fft_fft_SDFChainRadix22__GEN_1116); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1119 = 8'h1b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3c85) : $signed(fft_fft_SDFChainRadix22__GEN_1117); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1120 = 8'h1b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh14d2) : $signed(fft_fft_SDFChainRadix22__GEN_1118); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1121 = 8'h1c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_1119); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1122 = 8'h1c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_1120); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1123 = 8'h1d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3bfd) : $signed(fft_fft_SDFChainRadix22__GEN_1121); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1124 = 8'h1d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh164c) : $signed(fft_fft_SDFChainRadix22__GEN_1122); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1125 = 8'h1e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3bb6) : $signed(fft_fft_SDFChainRadix22__GEN_1123); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1126 = 8'h1e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1709) : $signed(fft_fft_SDFChainRadix22__GEN_1124); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1127 = 8'h1f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3b6d) : $signed(fft_fft_SDFChainRadix22__GEN_1125); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1128 = 8'h1f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh17c4) : $signed(fft_fft_SDFChainRadix22__GEN_1126); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1129 = 8'h20 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_1127); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1130 = 8'h20 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_1128); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1131 = 8'h21 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ad3) : $signed(fft_fft_SDFChainRadix22__GEN_1129); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1132 = 8'h21 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1937) : $signed(fft_fft_SDFChainRadix22__GEN_1130); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1133 = 8'h22 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3a82) : $signed(fft_fft_SDFChainRadix22__GEN_1131); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1134 = 8'h22 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh19ef) : $signed(fft_fft_SDFChainRadix22__GEN_1132); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1135 = 8'h23 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3a30) : $signed(fft_fft_SDFChainRadix22__GEN_1133); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1136 = 8'h23 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1aa7) : $signed(fft_fft_SDFChainRadix22__GEN_1134); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1137 = 8'h24 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_1135); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1138 = 8'h24 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_1136); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1139 = 8'h25 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3984) : $signed(fft_fft_SDFChainRadix22__GEN_1137); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1140 = 8'h25 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1c12) : $signed(fft_fft_SDFChainRadix22__GEN_1138); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1141 = 8'h26 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh392b) : $signed(fft_fft_SDFChainRadix22__GEN_1139); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1142 = 8'h26 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1cc6) : $signed(fft_fft_SDFChainRadix22__GEN_1140); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1143 = 8'h27 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh38cf) : $signed(fft_fft_SDFChainRadix22__GEN_1141); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1144 = 8'h27 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1d79) : $signed(fft_fft_SDFChainRadix22__GEN_1142); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1145 = 8'h28 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_1143); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1146 = 8'h28 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_1144); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1147 = 8'h29 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3812) : $signed(fft_fft_SDFChainRadix22__GEN_1145); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1148 = 8'h29 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1edc) : $signed(fft_fft_SDFChainRadix22__GEN_1146); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1149 = 8'h2a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh37b0) : $signed(fft_fft_SDFChainRadix22__GEN_1147); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1150 = 8'h2a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1f8c) : $signed(fft_fft_SDFChainRadix22__GEN_1148); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1151 = 8'h2b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh374b) : $signed(fft_fft_SDFChainRadix22__GEN_1149); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1152 = 8'h2b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh203a) : $signed(fft_fft_SDFChainRadix22__GEN_1150); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1153 = 8'h2c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_1151); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1154 = 8'h2c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_1152); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1155 = 8'h2d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh367d) : $signed(fft_fft_SDFChainRadix22__GEN_1153); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1156 = 8'h2d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2193) : $signed(fft_fft_SDFChainRadix22__GEN_1154); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1157 = 8'h2e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3612) : $signed(fft_fft_SDFChainRadix22__GEN_1155); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1158 = 8'h2e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh223d) : $signed(fft_fft_SDFChainRadix22__GEN_1156); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1159 = 8'h2f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh35a5) : $signed(fft_fft_SDFChainRadix22__GEN_1157); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1160 = 8'h2f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh22e7) : $signed(fft_fft_SDFChainRadix22__GEN_1158); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1161 = 8'h30 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_1159); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1162 = 8'h30 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_1160); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1163 = 8'h31 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh34c6) : $signed(fft_fft_SDFChainRadix22__GEN_1161); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1164 = 8'h31 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2435) : $signed(fft_fft_SDFChainRadix22__GEN_1162); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1165 = 8'h32 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3453) : $signed(fft_fft_SDFChainRadix22__GEN_1163); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1166 = 8'h32 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh24da) : $signed(fft_fft_SDFChainRadix22__GEN_1164); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1167 = 8'h33 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh33df) : $signed(fft_fft_SDFChainRadix22__GEN_1165); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1168 = 8'h33 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh257e) : $signed(fft_fft_SDFChainRadix22__GEN_1166); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1169 = 8'h34 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_1167); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1170 = 8'h34 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_1168); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1171 = 8'h35 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh32ef) : $signed(fft_fft_SDFChainRadix22__GEN_1169); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1172 = 8'h35 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh26c1) : $signed(fft_fft_SDFChainRadix22__GEN_1170); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1173 = 8'h36 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3274) : $signed(fft_fft_SDFChainRadix22__GEN_1171); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1174 = 8'h36 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2760) : $signed(fft_fft_SDFChainRadix22__GEN_1172); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1175 = 8'h37 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh31f8) : $signed(fft_fft_SDFChainRadix22__GEN_1173); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1176 = 8'h37 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh27fe) : $signed(fft_fft_SDFChainRadix22__GEN_1174); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1177 = 8'h38 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_1175); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1178 = 8'h38 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_1176); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1179 = 8'h39 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh30f9) : $signed(fft_fft_SDFChainRadix22__GEN_1177); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1180 = 8'h39 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2935) : $signed(fft_fft_SDFChainRadix22__GEN_1178); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1181 = 8'h3a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3076) : $signed(fft_fft_SDFChainRadix22__GEN_1179); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1182 = 8'h3a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh29ce) : $signed(fft_fft_SDFChainRadix22__GEN_1180); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1183 = 8'h3b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2ff2) : $signed(fft_fft_SDFChainRadix22__GEN_1181); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1184 = 8'h3b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2a65) : $signed(fft_fft_SDFChainRadix22__GEN_1182); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1185 = 8'h3c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_1183); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1186 = 8'h3c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_1184); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1187 = 8'h3d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2ee4) : $signed(fft_fft_SDFChainRadix22__GEN_1185); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1188 = 8'h3d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2b8f) : $signed(fft_fft_SDFChainRadix22__GEN_1186); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1189 = 8'h3e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2e5a) : $signed(fft_fft_SDFChainRadix22__GEN_1187); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1190 = 8'h3e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2c21) : $signed(fft_fft_SDFChainRadix22__GEN_1188); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1191 = 8'h3f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2dcf) : $signed(fft_fft_SDFChainRadix22__GEN_1189); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1192 = 8'h3f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2cb2) : $signed(fft_fft_SDFChainRadix22__GEN_1190); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1193 = 8'h40 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_1191); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1194 = 8'h40 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_1192); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1195 = 8'h41 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2cb2) : $signed(fft_fft_SDFChainRadix22__GEN_1193); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1196 = 8'h41 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2dcf) : $signed(fft_fft_SDFChainRadix22__GEN_1194); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1197 = 8'h42 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2c21) : $signed(fft_fft_SDFChainRadix22__GEN_1195); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1198 = 8'h42 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2e5a) : $signed(fft_fft_SDFChainRadix22__GEN_1196); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1199 = 8'h43 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2b8f) : $signed(fft_fft_SDFChainRadix22__GEN_1197); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1200 = 8'h43 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2ee4) : $signed(fft_fft_SDFChainRadix22__GEN_1198); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1201 = 8'h44 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_1199); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1202 = 8'h44 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_1200); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1203 = 8'h45 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2a65) : $signed(fft_fft_SDFChainRadix22__GEN_1201); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1204 = 8'h45 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2ff2) : $signed(fft_fft_SDFChainRadix22__GEN_1202); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1205 = 8'h46 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh29ce) : $signed(fft_fft_SDFChainRadix22__GEN_1203); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1206 = 8'h46 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3076) : $signed(fft_fft_SDFChainRadix22__GEN_1204); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1207 = 8'h47 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2935) : $signed(fft_fft_SDFChainRadix22__GEN_1205); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1208 = 8'h47 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh30f9) : $signed(fft_fft_SDFChainRadix22__GEN_1206); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1209 = 8'h48 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_1207); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1210 = 8'h48 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_1208); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1211 = 8'h49 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh27fe) : $signed(fft_fft_SDFChainRadix22__GEN_1209); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1212 = 8'h49 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh31f8) : $signed(fft_fft_SDFChainRadix22__GEN_1210); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1213 = 8'h4a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2760) : $signed(fft_fft_SDFChainRadix22__GEN_1211); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1214 = 8'h4a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3274) : $signed(fft_fft_SDFChainRadix22__GEN_1212); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1215 = 8'h4b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh26c1) : $signed(fft_fft_SDFChainRadix22__GEN_1213); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1216 = 8'h4b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh32ef) : $signed(fft_fft_SDFChainRadix22__GEN_1214); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1217 = 8'h4c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_1215); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1218 = 8'h4c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_1216); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1219 = 8'h4d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh257e) : $signed(fft_fft_SDFChainRadix22__GEN_1217); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1220 = 8'h4d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh33df) : $signed(fft_fft_SDFChainRadix22__GEN_1218); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1221 = 8'h4e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh24da) : $signed(fft_fft_SDFChainRadix22__GEN_1219); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1222 = 8'h4e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3453) : $signed(fft_fft_SDFChainRadix22__GEN_1220); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1223 = 8'h4f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2435) : $signed(fft_fft_SDFChainRadix22__GEN_1221); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1224 = 8'h4f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh34c6) : $signed(fft_fft_SDFChainRadix22__GEN_1222); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1225 = 8'h50 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_1223); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1226 = 8'h50 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_1224); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1227 = 8'h51 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh22e7) : $signed(fft_fft_SDFChainRadix22__GEN_1225); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1228 = 8'h51 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh35a5) : $signed(fft_fft_SDFChainRadix22__GEN_1226); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1229 = 8'h52 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh223d) : $signed(fft_fft_SDFChainRadix22__GEN_1227); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1230 = 8'h52 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3612) : $signed(fft_fft_SDFChainRadix22__GEN_1228); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1231 = 8'h53 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2193) : $signed(fft_fft_SDFChainRadix22__GEN_1229); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1232 = 8'h53 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh367d) : $signed(fft_fft_SDFChainRadix22__GEN_1230); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1233 = 8'h54 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_1231); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1234 = 8'h54 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_1232); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1235 = 8'h55 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh203a) : $signed(fft_fft_SDFChainRadix22__GEN_1233); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1236 = 8'h55 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh374b) : $signed(fft_fft_SDFChainRadix22__GEN_1234); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1237 = 8'h56 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1f8c) : $signed(fft_fft_SDFChainRadix22__GEN_1235); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1238 = 8'h56 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh37b0) : $signed(fft_fft_SDFChainRadix22__GEN_1236); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1239 = 8'h57 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1edc) : $signed(fft_fft_SDFChainRadix22__GEN_1237); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1240 = 8'h57 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3812) : $signed(fft_fft_SDFChainRadix22__GEN_1238); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1241 = 8'h58 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_1239); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1242 = 8'h58 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_1240); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1243 = 8'h59 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1d79) : $signed(fft_fft_SDFChainRadix22__GEN_1241); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1244 = 8'h59 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh38cf) : $signed(fft_fft_SDFChainRadix22__GEN_1242); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1245 = 8'h5a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1cc6) : $signed(fft_fft_SDFChainRadix22__GEN_1243); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1246 = 8'h5a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh392b) : $signed(fft_fft_SDFChainRadix22__GEN_1244); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1247 = 8'h5b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1c12) : $signed(fft_fft_SDFChainRadix22__GEN_1245); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1248 = 8'h5b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3984) : $signed(fft_fft_SDFChainRadix22__GEN_1246); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1249 = 8'h5c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_1247); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1250 = 8'h5c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_1248); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1251 = 8'h5d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1aa7) : $signed(fft_fft_SDFChainRadix22__GEN_1249); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1252 = 8'h5d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3a30) : $signed(fft_fft_SDFChainRadix22__GEN_1250); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1253 = 8'h5e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh19ef) : $signed(fft_fft_SDFChainRadix22__GEN_1251); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1254 = 8'h5e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3a82) : $signed(fft_fft_SDFChainRadix22__GEN_1252); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1255 = 8'h5f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1937) : $signed(fft_fft_SDFChainRadix22__GEN_1253); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1256 = 8'h5f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ad3) : $signed(fft_fft_SDFChainRadix22__GEN_1254); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1257 = 8'h60 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_1255); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1258 = 8'h60 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_1256); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1259 = 8'h61 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh17c4) : $signed(fft_fft_SDFChainRadix22__GEN_1257); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1260 = 8'h61 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3b6d) : $signed(fft_fft_SDFChainRadix22__GEN_1258); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1261 = 8'h62 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1709) : $signed(fft_fft_SDFChainRadix22__GEN_1259); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1262 = 8'h62 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3bb6) : $signed(fft_fft_SDFChainRadix22__GEN_1260); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1263 = 8'h63 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh164c) : $signed(fft_fft_SDFChainRadix22__GEN_1261); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1264 = 8'h63 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3bfd) : $signed(fft_fft_SDFChainRadix22__GEN_1262); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1265 = 8'h64 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_1263); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1266 = 8'h64 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_1264); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1267 = 8'h65 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh14d2) : $signed(fft_fft_SDFChainRadix22__GEN_1265); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1268 = 8'h65 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3c85) : $signed(fft_fft_SDFChainRadix22__GEN_1266); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1269 = 8'h66 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1413) : $signed(fft_fft_SDFChainRadix22__GEN_1267); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1270 = 8'h66 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3cc5) : $signed(fft_fft_SDFChainRadix22__GEN_1268); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1271 = 8'h67 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1354) : $signed(fft_fft_SDFChainRadix22__GEN_1269); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1272 = 8'h67 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d03) : $signed(fft_fft_SDFChainRadix22__GEN_1270); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1273 = 8'h68 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_1271); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1274 = 8'h68 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_1272); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1275 = 8'h69 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh11d3) : $signed(fft_fft_SDFChainRadix22__GEN_1273); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1276 = 8'h69 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d78) : $signed(fft_fft_SDFChainRadix22__GEN_1274); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1277 = 8'h6a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1112) : $signed(fft_fft_SDFChainRadix22__GEN_1275); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1278 = 8'h6a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3daf) : $signed(fft_fft_SDFChainRadix22__GEN_1276); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1279 = 8'h6b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1050) : $signed(fft_fft_SDFChainRadix22__GEN_1277); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1280 = 8'h6b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3de3) : $signed(fft_fft_SDFChainRadix22__GEN_1278); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1281 = 8'h6c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_1279); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1282 = 8'h6c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_1280); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1283 = 8'h6d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sheca) : $signed(fft_fft_SDFChainRadix22__GEN_1281); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1284 = 8'h6d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e45) : $signed(fft_fft_SDFChainRadix22__GEN_1282); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1285 = 8'h6e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'she06) : $signed(fft_fft_SDFChainRadix22__GEN_1283); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1286 = 8'h6e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e72) : $signed(fft_fft_SDFChainRadix22__GEN_1284); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1287 = 8'h6f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shd41) : $signed(fft_fft_SDFChainRadix22__GEN_1285); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1288 = 8'h6f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e9d) : $signed(fft_fft_SDFChainRadix22__GEN_1286); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1289 = 8'h70 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_1287); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1290 = 8'h70 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_1288); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1291 = 8'h71 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shbb7) : $signed(fft_fft_SDFChainRadix22__GEN_1289); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1292 = 8'h71 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3eeb) : $signed(fft_fft_SDFChainRadix22__GEN_1290); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1293 = 8'h72 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shaf1) : $signed(fft_fft_SDFChainRadix22__GEN_1291); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1294 = 8'h72 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f0f) : $signed(fft_fft_SDFChainRadix22__GEN_1292); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1295 = 8'h73 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sha2b) : $signed(fft_fft_SDFChainRadix22__GEN_1293); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1296 = 8'h73 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f30) : $signed(fft_fft_SDFChainRadix22__GEN_1294); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1297 = 8'h74 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_1295); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1298 = 8'h74 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_1296); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1299 = 8'h75 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh89d) : $signed(fft_fft_SDFChainRadix22__GEN_1297); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1300 = 8'h75 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f6b) : $signed(fft_fft_SDFChainRadix22__GEN_1298); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1301 = 8'h76 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh7d6) : $signed(fft_fft_SDFChainRadix22__GEN_1299); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1302 = 8'h76 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f85) : $signed(fft_fft_SDFChainRadix22__GEN_1300); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1303 = 8'h77 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh70e) : $signed(fft_fft_SDFChainRadix22__GEN_1301); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1304 = 8'h77 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f9c) : $signed(fft_fft_SDFChainRadix22__GEN_1302); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1305 = 8'h78 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_1303); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1306 = 8'h78 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_1304); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1307 = 8'h79 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh57e) : $signed(fft_fft_SDFChainRadix22__GEN_1305); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1308 = 8'h79 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fc4) : $signed(fft_fft_SDFChainRadix22__GEN_1306); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1309 = 8'h7a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh4b5) : $signed(fft_fft_SDFChainRadix22__GEN_1307); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1310 = 8'h7a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fd4) : $signed(fft_fft_SDFChainRadix22__GEN_1308); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1311 = 8'h7b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ed) : $signed(fft_fft_SDFChainRadix22__GEN_1309); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1312 = 8'h7b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fe1) : $signed(fft_fft_SDFChainRadix22__GEN_1310); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1313 = 8'h7c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh324) : $signed(fft_fft_SDFChainRadix22__GEN_1311); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1314 = 8'h7c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fec) : $signed(fft_fft_SDFChainRadix22__GEN_1312); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1315 = 8'h7d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh25b) : $signed(fft_fft_SDFChainRadix22__GEN_1313); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1316 = 8'h7d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ff5) : $signed(fft_fft_SDFChainRadix22__GEN_1314); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1317 = 8'h7e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh192) : $signed(fft_fft_SDFChainRadix22__GEN_1315); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1318 = 8'h7e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ffb) : $signed(fft_fft_SDFChainRadix22__GEN_1316); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1319 = 8'h7f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shc9) : $signed(fft_fft_SDFChainRadix22__GEN_1317); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1320 = 8'h7f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fff) : $signed(fft_fft_SDFChainRadix22__GEN_1318); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1321 = 8'h80 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh0) : $signed(fft_fft_SDFChainRadix22__GEN_1319); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1322 = 8'h80 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh4000) : $signed(fft_fft_SDFChainRadix22__GEN_1320); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1323 = 8'h81 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shc9) : $signed(fft_fft_SDFChainRadix22__GEN_1321); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1324 = 8'h81 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fff) : $signed(fft_fft_SDFChainRadix22__GEN_1322); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1325 = 8'h82 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh192) : $signed(fft_fft_SDFChainRadix22__GEN_1323); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1326 = 8'h82 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ffb) : $signed(fft_fft_SDFChainRadix22__GEN_1324); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1327 = 8'h83 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh324) : $signed(fft_fft_SDFChainRadix22__GEN_1325); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1328 = 8'h83 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fec) : $signed(fft_fft_SDFChainRadix22__GEN_1326); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1329 = 8'h84 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh4b5) : $signed(fft_fft_SDFChainRadix22__GEN_1327); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1330 = 8'h84 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fd4) : $signed(fft_fft_SDFChainRadix22__GEN_1328); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1331 = 8'h85 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh57e) : $signed(fft_fft_SDFChainRadix22__GEN_1329); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1332 = 8'h85 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fc4) : $signed(fft_fft_SDFChainRadix22__GEN_1330); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1333 = 8'h86 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_1331); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1334 = 8'h86 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_1332); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1335 = 8'h87 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh7d6) : $signed(fft_fft_SDFChainRadix22__GEN_1333); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1336 = 8'h87 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f85) : $signed(fft_fft_SDFChainRadix22__GEN_1334); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1337 = 8'h88 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_1335); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1338 = 8'h88 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_1336); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1339 = 8'h89 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sha2b) : $signed(fft_fft_SDFChainRadix22__GEN_1337); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1340 = 8'h89 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f30) : $signed(fft_fft_SDFChainRadix22__GEN_1338); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1341 = 8'h8a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shaf1) : $signed(fft_fft_SDFChainRadix22__GEN_1339); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1342 = 8'h8a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f0f) : $signed(fft_fft_SDFChainRadix22__GEN_1340); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1343 = 8'h8b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_1341); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1344 = 8'h8b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_1342); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1345 = 8'h8c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'she06) : $signed(fft_fft_SDFChainRadix22__GEN_1343); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1346 = 8'h8c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e72) : $signed(fft_fft_SDFChainRadix22__GEN_1344); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1347 = 8'h8d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sheca) : $signed(fft_fft_SDFChainRadix22__GEN_1345); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1348 = 8'h8d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e45) : $signed(fft_fft_SDFChainRadix22__GEN_1346); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1349 = 8'h8e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_1347); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1350 = 8'h8e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_1348); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1351 = 8'h8f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1112) : $signed(fft_fft_SDFChainRadix22__GEN_1349); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1352 = 8'h8f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3daf) : $signed(fft_fft_SDFChainRadix22__GEN_1350); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1353 = 8'h90 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_1351); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1354 = 8'h90 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_1352); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1355 = 8'h91 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1354) : $signed(fft_fft_SDFChainRadix22__GEN_1353); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1356 = 8'h91 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d03) : $signed(fft_fft_SDFChainRadix22__GEN_1354); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1357 = 8'h92 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1413) : $signed(fft_fft_SDFChainRadix22__GEN_1355); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1358 = 8'h92 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3cc5) : $signed(fft_fft_SDFChainRadix22__GEN_1356); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1359 = 8'h93 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_1357); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1360 = 8'h93 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_1358); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1361 = 8'h94 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1709) : $signed(fft_fft_SDFChainRadix22__GEN_1359); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1362 = 8'h94 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3bb6) : $signed(fft_fft_SDFChainRadix22__GEN_1360); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1363 = 8'h95 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh17c4) : $signed(fft_fft_SDFChainRadix22__GEN_1361); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1364 = 8'h95 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3b6d) : $signed(fft_fft_SDFChainRadix22__GEN_1362); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1365 = 8'h96 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_1363); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1366 = 8'h96 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_1364); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1367 = 8'h97 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh19ef) : $signed(fft_fft_SDFChainRadix22__GEN_1365); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1368 = 8'h97 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3a82) : $signed(fft_fft_SDFChainRadix22__GEN_1366); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1369 = 8'h98 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_1367); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1370 = 8'h98 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_1368); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1371 = 8'h99 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1c12) : $signed(fft_fft_SDFChainRadix22__GEN_1369); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1372 = 8'h99 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3984) : $signed(fft_fft_SDFChainRadix22__GEN_1370); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1373 = 8'h9a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1cc6) : $signed(fft_fft_SDFChainRadix22__GEN_1371); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1374 = 8'h9a == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh392b) : $signed(fft_fft_SDFChainRadix22__GEN_1372); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1375 = 8'h9b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_1373); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1376 = 8'h9b == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_1374); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1377 = 8'h9c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1f8c) : $signed(fft_fft_SDFChainRadix22__GEN_1375); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1378 = 8'h9c == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh37b0) : $signed(fft_fft_SDFChainRadix22__GEN_1376); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1379 = 8'h9d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh203a) : $signed(fft_fft_SDFChainRadix22__GEN_1377); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1380 = 8'h9d == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh374b) : $signed(fft_fft_SDFChainRadix22__GEN_1378); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1381 = 8'h9e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_1379); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1382 = 8'h9e == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_1380); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1383 = 8'h9f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh223d) : $signed(fft_fft_SDFChainRadix22__GEN_1381); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1384 = 8'h9f == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3612) : $signed(fft_fft_SDFChainRadix22__GEN_1382); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1385 = 8'ha0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_1383); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1386 = 8'ha0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_1384); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1387 = 8'ha1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2435) : $signed(fft_fft_SDFChainRadix22__GEN_1385); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1388 = 8'ha1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh34c6) : $signed(fft_fft_SDFChainRadix22__GEN_1386); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1389 = 8'ha2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh24da) : $signed(fft_fft_SDFChainRadix22__GEN_1387); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1390 = 8'ha2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3453) : $signed(fft_fft_SDFChainRadix22__GEN_1388); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1391 = 8'ha3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_1389); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1392 = 8'ha3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_1390); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1393 = 8'ha4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2760) : $signed(fft_fft_SDFChainRadix22__GEN_1391); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1394 = 8'ha4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3274) : $signed(fft_fft_SDFChainRadix22__GEN_1392); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1395 = 8'ha5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh27fe) : $signed(fft_fft_SDFChainRadix22__GEN_1393); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1396 = 8'ha5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh31f8) : $signed(fft_fft_SDFChainRadix22__GEN_1394); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1397 = 8'ha6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_1395); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1398 = 8'ha6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_1396); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1399 = 8'ha7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh29ce) : $signed(fft_fft_SDFChainRadix22__GEN_1397); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1400 = 8'ha7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3076) : $signed(fft_fft_SDFChainRadix22__GEN_1398); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1401 = 8'ha8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_1399); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1402 = 8'ha8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_1400); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1403 = 8'ha9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2b8f) : $signed(fft_fft_SDFChainRadix22__GEN_1401); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1404 = 8'ha9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2ee4) : $signed(fft_fft_SDFChainRadix22__GEN_1402); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1405 = 8'haa == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2c21) : $signed(fft_fft_SDFChainRadix22__GEN_1403); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1406 = 8'haa == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2e5a) : $signed(fft_fft_SDFChainRadix22__GEN_1404); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1407 = 8'hab == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_1405); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1408 = 8'hab == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2d41) : $signed(fft_fft_SDFChainRadix22__GEN_1406); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1409 = 8'hac == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2e5a) : $signed(fft_fft_SDFChainRadix22__GEN_1407); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1410 = 8'hac == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2c21) : $signed(fft_fft_SDFChainRadix22__GEN_1408); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1411 = 8'had == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2ee4) : $signed(fft_fft_SDFChainRadix22__GEN_1409); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1412 = 8'had == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2b8f) : $signed(fft_fft_SDFChainRadix22__GEN_1410); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1413 = 8'hae == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_1411); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1414 = 8'hae == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_1412); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1415 = 8'haf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3076) : $signed(fft_fft_SDFChainRadix22__GEN_1413); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1416 = 8'haf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh29ce) : $signed(fft_fft_SDFChainRadix22__GEN_1414); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1417 = 8'hb0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_1415); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1418 = 8'hb0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_1416); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1419 = 8'hb1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh31f8) : $signed(fft_fft_SDFChainRadix22__GEN_1417); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1420 = 8'hb1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh27fe) : $signed(fft_fft_SDFChainRadix22__GEN_1418); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1421 = 8'hb2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3274) : $signed(fft_fft_SDFChainRadix22__GEN_1419); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1422 = 8'hb2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2760) : $signed(fft_fft_SDFChainRadix22__GEN_1420); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1423 = 8'hb3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3368) : $signed(fft_fft_SDFChainRadix22__GEN_1421); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1424 = 8'hb3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2620) : $signed(fft_fft_SDFChainRadix22__GEN_1422); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1425 = 8'hb4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3453) : $signed(fft_fft_SDFChainRadix22__GEN_1423); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1426 = 8'hb4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh24da) : $signed(fft_fft_SDFChainRadix22__GEN_1424); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1427 = 8'hb5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh34c6) : $signed(fft_fft_SDFChainRadix22__GEN_1425); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1428 = 8'hb5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2435) : $signed(fft_fft_SDFChainRadix22__GEN_1426); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1429 = 8'hb6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_1427); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1430 = 8'hb6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_1428); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1431 = 8'hb7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3612) : $signed(fft_fft_SDFChainRadix22__GEN_1429); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1432 = 8'hb7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh223d) : $signed(fft_fft_SDFChainRadix22__GEN_1430); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1433 = 8'hb8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_1431); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1434 = 8'hb8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_1432); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1435 = 8'hb9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh374b) : $signed(fft_fft_SDFChainRadix22__GEN_1433); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1436 = 8'hb9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh203a) : $signed(fft_fft_SDFChainRadix22__GEN_1434); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1437 = 8'hba == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh37b0) : $signed(fft_fft_SDFChainRadix22__GEN_1435); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1438 = 8'hba == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1f8c) : $signed(fft_fft_SDFChainRadix22__GEN_1436); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1439 = 8'hbb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3871) : $signed(fft_fft_SDFChainRadix22__GEN_1437); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1440 = 8'hbb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1e2b) : $signed(fft_fft_SDFChainRadix22__GEN_1438); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1441 = 8'hbc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh392b) : $signed(fft_fft_SDFChainRadix22__GEN_1439); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1442 = 8'hbc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1cc6) : $signed(fft_fft_SDFChainRadix22__GEN_1440); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1443 = 8'hbd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3984) : $signed(fft_fft_SDFChainRadix22__GEN_1441); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1444 = 8'hbd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1c12) : $signed(fft_fft_SDFChainRadix22__GEN_1442); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1445 = 8'hbe == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_1443); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1446 = 8'hbe == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_1444); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1447 = 8'hbf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3a82) : $signed(fft_fft_SDFChainRadix22__GEN_1445); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1448 = 8'hbf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh19ef) : $signed(fft_fft_SDFChainRadix22__GEN_1446); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1449 = 8'hc0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_1447); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1450 = 8'hc0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_1448); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1451 = 8'hc1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3b6d) : $signed(fft_fft_SDFChainRadix22__GEN_1449); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1452 = 8'hc1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh17c4) : $signed(fft_fft_SDFChainRadix22__GEN_1450); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1453 = 8'hc2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3bb6) : $signed(fft_fft_SDFChainRadix22__GEN_1451); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1454 = 8'hc2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1709) : $signed(fft_fft_SDFChainRadix22__GEN_1452); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1455 = 8'hc3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3c42) : $signed(fft_fft_SDFChainRadix22__GEN_1453); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1456 = 8'hc3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1590) : $signed(fft_fft_SDFChainRadix22__GEN_1454); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1457 = 8'hc4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3cc5) : $signed(fft_fft_SDFChainRadix22__GEN_1455); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1458 = 8'hc4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1413) : $signed(fft_fft_SDFChainRadix22__GEN_1456); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1459 = 8'hc5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d03) : $signed(fft_fft_SDFChainRadix22__GEN_1457); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1460 = 8'hc5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1354) : $signed(fft_fft_SDFChainRadix22__GEN_1458); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1461 = 8'hc6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_1459); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1462 = 8'hc6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_1460); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1463 = 8'hc7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3daf) : $signed(fft_fft_SDFChainRadix22__GEN_1461); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1464 = 8'hc7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1112) : $signed(fft_fft_SDFChainRadix22__GEN_1462); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1465 = 8'hc8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_1463); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1466 = 8'hc8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_1464); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1467 = 8'hc9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e45) : $signed(fft_fft_SDFChainRadix22__GEN_1465); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1468 = 8'hc9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sheca) : $signed(fft_fft_SDFChainRadix22__GEN_1466); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1469 = 8'hca == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e72) : $signed(fft_fft_SDFChainRadix22__GEN_1467); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1470 = 8'hca == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'she06) : $signed(fft_fft_SDFChainRadix22__GEN_1468); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1471 = 8'hcb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ec5) : $signed(fft_fft_SDFChainRadix22__GEN_1469); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1472 = 8'hcb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shc7c) : $signed(fft_fft_SDFChainRadix22__GEN_1470); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1473 = 8'hcc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f0f) : $signed(fft_fft_SDFChainRadix22__GEN_1471); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1474 = 8'hcc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shaf1) : $signed(fft_fft_SDFChainRadix22__GEN_1472); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1475 = 8'hcd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f30) : $signed(fft_fft_SDFChainRadix22__GEN_1473); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1476 = 8'hcd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sha2b) : $signed(fft_fft_SDFChainRadix22__GEN_1474); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1477 = 8'hce == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_1475); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1478 = 8'hce == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_1476); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1479 = 8'hcf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f85) : $signed(fft_fft_SDFChainRadix22__GEN_1477); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1480 = 8'hcf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh7d6) : $signed(fft_fft_SDFChainRadix22__GEN_1478); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1481 = 8'hd0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_1479); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1482 = 8'hd0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_1480); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1483 = 8'hd1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fc4) : $signed(fft_fft_SDFChainRadix22__GEN_1481); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1484 = 8'hd1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh57e) : $signed(fft_fft_SDFChainRadix22__GEN_1482); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1485 = 8'hd2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fd4) : $signed(fft_fft_SDFChainRadix22__GEN_1483); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1486 = 8'hd2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh4b5) : $signed(fft_fft_SDFChainRadix22__GEN_1484); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1487 = 8'hd3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fec) : $signed(fft_fft_SDFChainRadix22__GEN_1485); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1488 = 8'hd3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh324) : $signed(fft_fft_SDFChainRadix22__GEN_1486); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1489 = 8'hd4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ffb) : $signed(fft_fft_SDFChainRadix22__GEN_1487); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1490 = 8'hd4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh192) : $signed(fft_fft_SDFChainRadix22__GEN_1488); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1491 = 8'hd5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fff) : $signed(fft_fft_SDFChainRadix22__GEN_1489); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1492 = 8'hd5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shc9) : $signed(fft_fft_SDFChainRadix22__GEN_1490); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1493 = 8'hd6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3ffb) : $signed(fft_fft_SDFChainRadix22__GEN_1491); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1494 = 8'hd6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh192) : $signed(fft_fft_SDFChainRadix22__GEN_1492); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1495 = 8'hd7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fe1) : $signed(fft_fft_SDFChainRadix22__GEN_1493); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1496 = 8'hd7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ed) : $signed(fft_fft_SDFChainRadix22__GEN_1494); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1497 = 8'hd8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3fb1) : $signed(fft_fft_SDFChainRadix22__GEN_1495); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1498 = 8'hd8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh646) : $signed(fft_fft_SDFChainRadix22__GEN_1496); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1499 = 8'hd9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f6b) : $signed(fft_fft_SDFChainRadix22__GEN_1497); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1500 = 8'hd9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh89d) : $signed(fft_fft_SDFChainRadix22__GEN_1498); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1501 = 8'hda == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3f0f) : $signed(fft_fft_SDFChainRadix22__GEN_1499); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1502 = 8'hda == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shaf1) : $signed(fft_fft_SDFChainRadix22__GEN_1500); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1503 = 8'hdb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e9d) : $signed(fft_fft_SDFChainRadix22__GEN_1501); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1504 = 8'hdb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shd41) : $signed(fft_fft_SDFChainRadix22__GEN_1502); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1505 = 8'hdc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3e15) : $signed(fft_fft_SDFChainRadix22__GEN_1503); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1506 = 8'hdc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'shf8d) : $signed(fft_fft_SDFChainRadix22__GEN_1504); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1507 = 8'hdd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3d78) : $signed(fft_fft_SDFChainRadix22__GEN_1505); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1508 = 8'hdd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh11d3) : $signed(fft_fft_SDFChainRadix22__GEN_1506); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1509 = 8'hde == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3cc5) : $signed(fft_fft_SDFChainRadix22__GEN_1507); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1510 = 8'hde == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1413) : $signed(fft_fft_SDFChainRadix22__GEN_1508); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1511 = 8'hdf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3bfd) : $signed(fft_fft_SDFChainRadix22__GEN_1509); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1512 = 8'hdf == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh164c) : $signed(fft_fft_SDFChainRadix22__GEN_1510); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1513 = 8'he0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3b21) : $signed(fft_fft_SDFChainRadix22__GEN_1511); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1514 = 8'he0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh187e) : $signed(fft_fft_SDFChainRadix22__GEN_1512); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1515 = 8'he1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3a30) : $signed(fft_fft_SDFChainRadix22__GEN_1513); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1516 = 8'he1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1aa7) : $signed(fft_fft_SDFChainRadix22__GEN_1514); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1517 = 8'he2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh392b) : $signed(fft_fft_SDFChainRadix22__GEN_1515); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1518 = 8'he2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1cc6) : $signed(fft_fft_SDFChainRadix22__GEN_1516); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1519 = 8'he3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3812) : $signed(fft_fft_SDFChainRadix22__GEN_1517); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1520 = 8'he3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh1edc) : $signed(fft_fft_SDFChainRadix22__GEN_1518); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1521 = 8'he4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh36e5) : $signed(fft_fft_SDFChainRadix22__GEN_1519); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1522 = 8'he4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh20e7) : $signed(fft_fft_SDFChainRadix22__GEN_1520); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1523 = 8'he5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh35a5) : $signed(fft_fft_SDFChainRadix22__GEN_1521); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1524 = 8'he5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh22e7) : $signed(fft_fft_SDFChainRadix22__GEN_1522); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1525 = 8'he6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3453) : $signed(fft_fft_SDFChainRadix22__GEN_1523); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1526 = 8'he6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh24da) : $signed(fft_fft_SDFChainRadix22__GEN_1524); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1527 = 8'he7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh32ef) : $signed(fft_fft_SDFChainRadix22__GEN_1525); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1528 = 8'he7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh26c1) : $signed(fft_fft_SDFChainRadix22__GEN_1526); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1529 = 8'he8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh3179) : $signed(fft_fft_SDFChainRadix22__GEN_1527); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1530 = 8'he8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh289a) : $signed(fft_fft_SDFChainRadix22__GEN_1528); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1531 = 8'he9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2ff2) : $signed(fft_fft_SDFChainRadix22__GEN_1529); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1532 = 8'he9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2a65) : $signed(fft_fft_SDFChainRadix22__GEN_1530); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1533 = 8'hea == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2e5a) : $signed(fft_fft_SDFChainRadix22__GEN_1531); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1534 = 8'hea == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2c21) : $signed(fft_fft_SDFChainRadix22__GEN_1532); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1535 = 8'heb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2cb2) : $signed(fft_fft_SDFChainRadix22__GEN_1533); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1536 = 8'heb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2dcf) : $signed(fft_fft_SDFChainRadix22__GEN_1534); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1537 = 8'hec == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2afb) : $signed(fft_fft_SDFChainRadix22__GEN_1535); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1538 = 8'hec == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh2f6c) : $signed(fft_fft_SDFChainRadix22__GEN_1536); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1539 = 8'hed == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2935) : $signed(fft_fft_SDFChainRadix22__GEN_1537); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1540 = 8'hed == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh30f9) : $signed(fft_fft_SDFChainRadix22__GEN_1538); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1541 = 8'hee == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2760) : $signed(fft_fft_SDFChainRadix22__GEN_1539); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1542 = 8'hee == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3274) : $signed(fft_fft_SDFChainRadix22__GEN_1540); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1543 = 8'hef == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh257e) : $signed(fft_fft_SDFChainRadix22__GEN_1541); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1544 = 8'hef == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh33df) : $signed(fft_fft_SDFChainRadix22__GEN_1542); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1545 = 8'hf0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh238e) : $signed(fft_fft_SDFChainRadix22__GEN_1543); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1546 = 8'hf0 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3537) : $signed(fft_fft_SDFChainRadix22__GEN_1544); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1547 = 8'hf1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh2193) : $signed(fft_fft_SDFChainRadix22__GEN_1545); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1548 = 8'hf1 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh367d) : $signed(fft_fft_SDFChainRadix22__GEN_1546); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1549 = 8'hf2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1f8c) : $signed(fft_fft_SDFChainRadix22__GEN_1547); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1550 = 8'hf2 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh37b0) : $signed(fft_fft_SDFChainRadix22__GEN_1548); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1551 = 8'hf3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1d79) : $signed(fft_fft_SDFChainRadix22__GEN_1549); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1552 = 8'hf3 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh38cf) : $signed(fft_fft_SDFChainRadix22__GEN_1550); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1553 = 8'hf4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1b5d) : $signed(fft_fft_SDFChainRadix22__GEN_1551); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1554 = 8'hf4 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh39db) : $signed(fft_fft_SDFChainRadix22__GEN_1552); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1555 = 8'hf5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1937) : $signed(fft_fft_SDFChainRadix22__GEN_1553); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1556 = 8'hf5 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ad3) : $signed(fft_fft_SDFChainRadix22__GEN_1554); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1557 = 8'hf6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1709) : $signed(fft_fft_SDFChainRadix22__GEN_1555); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1558 = 8'hf6 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3bb6) : $signed(fft_fft_SDFChainRadix22__GEN_1556); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1559 = 8'hf7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh14d2) : $signed(fft_fft_SDFChainRadix22__GEN_1557); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1560 = 8'hf7 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3c85) : $signed(fft_fft_SDFChainRadix22__GEN_1558); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1561 = 8'hf8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1294) : $signed(fft_fft_SDFChainRadix22__GEN_1559); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1562 = 8'hf8 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3d3f) : $signed(fft_fft_SDFChainRadix22__GEN_1560); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1563 = 8'hf9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh1050) : $signed(fft_fft_SDFChainRadix22__GEN_1561); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1564 = 8'hf9 == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3de3) : $signed(fft_fft_SDFChainRadix22__GEN_1562); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1565 = 8'hfa == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'she06) : $signed(fft_fft_SDFChainRadix22__GEN_1563); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1566 = 8'hfa == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3e72) : $signed(fft_fft_SDFChainRadix22__GEN_1564); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1567 = 8'hfb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'shbb7) : $signed(fft_fft_SDFChainRadix22__GEN_1565); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1568 = 8'hfb == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3eeb) : $signed(fft_fft_SDFChainRadix22__GEN_1566); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1569 = 8'hfc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh964) : $signed(fft_fft_SDFChainRadix22__GEN_1567); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1570 = 8'hfc == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f4f) : $signed(fft_fft_SDFChainRadix22__GEN_1568); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1571 = 8'hfd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh70e) : $signed(fft_fft_SDFChainRadix22__GEN_1569); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1572 = 8'hfd == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3f9c) : $signed(fft_fft_SDFChainRadix22__GEN_1570); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1573 = 8'hfe == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh4b5) : $signed(fft_fft_SDFChainRadix22__GEN_1571); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1574 = 8'hfe == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3fd4) : $signed(fft_fft_SDFChainRadix22__GEN_1572); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__GEN_1575 = 8'hff == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(-16'sh25b) : $signed(fft_fft_SDFChainRadix22__GEN_1573); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22_twiddles_7_imag = 8'hff == fft_fft_SDFChainRadix22__GEN_1064 ? $signed(16'sh3ff5) : $signed(fft_fft_SDFChainRadix22__GEN_1574); // @[SDFChainRadix22.scala 291:27]
  assign fft_fft_SDFChainRadix22__T_2096 = $signed(fft_fft_SDFChainRadix22__GEN_1575) + $signed(fft_fft_SDFChainRadix22_twiddles_7_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22_outputWires_6_real = fft_fft_SDFChainRadix22_sdf_stages_6_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22_outputWires_6_imag = fft_fft_SDFChainRadix22_sdf_stages_6_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22__T_2097 = $signed(fft_fft_SDFChainRadix22_outputWires_6_real) + $signed(fft_fft_SDFChainRadix22_outputWires_6_imag); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_2098 = $signed(fft_fft_SDFChainRadix22_outputWires_6_imag) - $signed(fft_fft_SDFChainRadix22_outputWires_6_real); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__GEN_2121 = {{1{fft_fft_SDFChainRadix22_outputWires_6_real[15]}},fft_fft_SDFChainRadix22_outputWires_6_real}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_2099 = $signed(fft_fft_SDFChainRadix22__GEN_2121) * $signed(fft_fft_SDFChainRadix22__T_2096); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2122 = {{1{fft_fft_SDFChainRadix22_twiddles_7_imag[15]}},fft_fft_SDFChainRadix22_twiddles_7_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_2100 = $signed(fft_fft_SDFChainRadix22__T_2097) * $signed(fft_fft_SDFChainRadix22__GEN_2122); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__GEN_2123 = {{1{fft_fft_SDFChainRadix22__GEN_1575[15]}},fft_fft_SDFChainRadix22__GEN_1575}; // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_2101 = $signed(fft_fft_SDFChainRadix22__T_2098) * $signed(fft_fft_SDFChainRadix22__GEN_2123); // @[FixedPointTypeClass.scala 211:35]
  assign fft_fft_SDFChainRadix22__T_2102 = $signed(fft_fft_SDFChainRadix22__T_2099) - $signed(fft_fft_SDFChainRadix22__T_2100); // @[FixedPointTypeClass.scala 33:22]
  assign fft_fft_SDFChainRadix22__T_2103 = $signed(fft_fft_SDFChainRadix22__T_2099) + $signed(fft_fft_SDFChainRadix22__T_2101); // @[FixedPointTypeClass.scala 24:22]
  assign fft_fft_SDFChainRadix22__T_2109 = $signed(fft_fft_SDFChainRadix22__T_2102) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_2110 = fft_fft_SDFChainRadix22__T_2109[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_2113 = $signed(fft_fft_SDFChainRadix22__T_2103) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign fft_fft_SDFChainRadix22__T_2114 = fft_fft_SDFChainRadix22__T_2113[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign fft_fft_SDFChainRadix22__T_2121 = fft_fft_SDFChainRadix22_sdf_stages_8_io_cntr < 9'h100; // @[SDFChainRadix22.scala 328:32]
  assign fft_fft_SDFChainRadix22__T_2122 = fft_fft_SDFChainRadix22_sdf_stages_8_io_cntr < 9'h180; // @[SDFChainRadix22.scala 328:78]
  assign fft_fft_SDFChainRadix22__T_2123 = fft_fft_SDFChainRadix22__T_2122 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign fft_fft_SDFChainRadix22__T_2124 = fft_fft_SDFChainRadix22__T_2121 ? 1'h0 : fft_fft_SDFChainRadix22__T_2123; // @[SDFChainRadix22.scala 328:19]
  assign fft_fft_SDFChainRadix22_outputWires_7_real = fft_fft_SDFChainRadix22_sdf_stages_7_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__T_2130 = 16'sh0 - $signed(fft_fft_SDFChainRadix22_outputWires_7_real); // @[FixedPointTypeClass.scala 39:43]
  assign fft_fft_SDFChainRadix22_outputWires_7_imag = fft_fft_SDFChainRadix22_sdf_stages_7_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign fft_fft_SDFChainRadix22__GEN_2091 = 4'h1 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_1_real) : $signed(fft_fft_SDFChainRadix22_outputWires_0_real); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2092 = 4'h1 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_1_imag) : $signed(fft_fft_SDFChainRadix22_outputWires_0_imag); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2093 = 4'h2 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_2_real) : $signed(fft_fft_SDFChainRadix22__GEN_2091); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2094 = 4'h2 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_2_imag) : $signed(fft_fft_SDFChainRadix22__GEN_2092); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2095 = 4'h3 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_3_real) : $signed(fft_fft_SDFChainRadix22__GEN_2093); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2096 = 4'h3 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_3_imag) : $signed(fft_fft_SDFChainRadix22__GEN_2094); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2097 = 4'h4 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_4_real) : $signed(fft_fft_SDFChainRadix22__GEN_2095); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2098 = 4'h4 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_4_imag) : $signed(fft_fft_SDFChainRadix22__GEN_2096); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2099 = 4'h5 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_5_real) : $signed(fft_fft_SDFChainRadix22__GEN_2097); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2100 = 4'h5 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_5_imag) : $signed(fft_fft_SDFChainRadix22__GEN_2098); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2101 = 4'h6 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_6_real) : $signed(fft_fft_SDFChainRadix22__GEN_2099); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2102 = 4'h6 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_6_imag) : $signed(fft_fft_SDFChainRadix22__GEN_2100); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2103 = 4'h7 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_7_real) : $signed(fft_fft_SDFChainRadix22__GEN_2101); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__GEN_2104 = 4'h7 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_7_imag) : $signed(fft_fft_SDFChainRadix22__GEN_2102); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22_outputWires_8_real = fft_fft_SDFChainRadix22_sdf_stages_8_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22__GEN_2105 = 4'h8 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_8_real) : $signed(fft_fft_SDFChainRadix22__GEN_2103); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22_outputWires_8_imag = fft_fft_SDFChainRadix22_sdf_stages_8_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign fft_fft_SDFChainRadix22__GEN_2106 = 4'h8 == fft_fft_SDFChainRadix22__T_49 ? $signed(fft_fft_SDFChainRadix22_outputWires_8_imag) : $signed(fft_fft_SDFChainRadix22__GEN_2104); // @[SDFChainRadix22.scala 364:24]
  assign fft_fft_SDFChainRadix22__T_2140 = ~fft_fft_SDFChainRadix22_initialOutDone; // @[SDFChainRadix22.scala 368:33]
  assign fft_fft_SDFChainRadix22__T_2141 = fft_fft_SDFChainRadix22_state != 2'h2; // @[SDFChainRadix22.scala 368:127]
  assign fft_fft_SDFChainRadix22__T_2142 = fft_fft_SDFChainRadix22_io_out_ready & fft_fft_SDFChainRadix22__T_2141; // @[SDFChainRadix22.scala 368:117]
  assign fft_fft_SDFChainRadix22__GEN_2124 = {$signed(fft_fft_SDFChainRadix22__GEN_2106), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  assign fft_fft_SDFChainRadix22__GEN_2107 = {{2{fft_fft_SDFChainRadix22__GEN_2124[29]}},fft_fft_SDFChainRadix22__GEN_2124}; // @[SDFChainRadix22.scala 375:33]
  assign fft_fft_SDFChainRadix22__GEN_2125 = {$signed(fft_fft_SDFChainRadix22__GEN_2105), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  assign fft_fft_SDFChainRadix22__GEN_2108 = {{2{fft_fft_SDFChainRadix22__GEN_2125[29]}},fft_fft_SDFChainRadix22__GEN_2125}; // @[SDFChainRadix22.scala 375:33]
  assign fft_fft_SDFChainRadix22__GEN_2126 = fft_fft_SDFChainRadix22__GEN_2108[31:14]; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 396:27]
  assign fft_fft_SDFChainRadix22__GEN_2128 = fft_fft_SDFChainRadix22__GEN_2107[31:14]; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 397:27]
  assign fft_fft_SDFChainRadix22_io_in_ready = fft_fft_SDFChainRadix22__T_2140 | fft_fft_SDFChainRadix22__T_2142; // @[SDFChainRadix22.scala 368:15]
  assign fft_fft_SDFChainRadix22_io_out_valid = fft_fft_SDFChainRadix22_enableInit & fft_fft_SDFChainRadix22_initialOutDone; // @[SDFChainRadix22.scala 401:18]
  assign fft_fft_SDFChainRadix22_io_out_bits_real = fft_fft_SDFChainRadix22__GEN_2126[15:0]; // @[SDFChainRadix22.scala 400:17]
  assign fft_fft_SDFChainRadix22_io_out_bits_imag = fft_fft_SDFChainRadix22__GEN_2128[15:0]; // @[SDFChainRadix22.scala 400:17]
  assign fft_fft_SDFChainRadix22_io_lastOut = fft_fft_SDFChainRadix22_pktEnd & fft_fft_SDFChainRadix22__T_83; // @[SDFChainRadix22.scala 428:14]
  assign fft_fft_SDFChainRadix22_io_busy = fft_fft_SDFChainRadix22_state != 2'h0; // @[SDFChainRadix22.scala 430:11]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_0_io_in_real = fft_fft_SDFChainRadix22_io_in_bits_real; // @[SDFChainRadix22.scala 347:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_io_in_imag = fft_fft_SDFChainRadix22_io_in_bits_imag; // @[SDFChainRadix22.scala 347:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_io_cntr = {{8'd0}, fft_fft_SDFChainRadix22__T_167}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_0_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_1_io_in_real = fft_fft_SDFChainRadix22__T_275[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_io_in_imag = fft_fft_SDFChainRadix22__T_279[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_io_cntr = {{7'd0}, fft_fft_SDFChainRadix22__T_174}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_1_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_2_io_in_real = fft_fft_SDFChainRadix22__T_289 ? $signed(fft_fft_SDFChainRadix22_outputWires_1_imag) : $signed(fft_fft_SDFChainRadix22_outputWires_1_real); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_io_in_imag = fft_fft_SDFChainRadix22__T_289 ? $signed(fft_fft_SDFChainRadix22__T_295) : $signed(fft_fft_SDFChainRadix22_outputWires_1_imag); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_io_cntr = {{6'd0}, fft_fft_SDFChainRadix22__T_181}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_2_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_3_io_in_real = fft_fft_SDFChainRadix22__T_407[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_io_in_imag = fft_fft_SDFChainRadix22__T_411[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_io_cntr = {{5'd0}, fft_fft_SDFChainRadix22__T_188}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_3_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_4_io_in_real = fft_fft_SDFChainRadix22__T_421 ? $signed(fft_fft_SDFChainRadix22_outputWires_3_imag) : $signed(fft_fft_SDFChainRadix22_outputWires_3_real); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_io_in_imag = fft_fft_SDFChainRadix22__T_421 ? $signed(fft_fft_SDFChainRadix22__T_427) : $signed(fft_fft_SDFChainRadix22_outputWires_3_imag); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_io_cntr = {{4'd0}, fft_fft_SDFChainRadix22__T_195}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_4_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_5_io_in_real = fft_fft_SDFChainRadix22__T_779[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_io_in_imag = fft_fft_SDFChainRadix22__T_783[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_io_cntr = {{3'd0}, fft_fft_SDFChainRadix22__T_202}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_5_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_6_io_in_real = fft_fft_SDFChainRadix22__T_793 ? $signed(fft_fft_SDFChainRadix22_outputWires_5_imag) : $signed(fft_fft_SDFChainRadix22_outputWires_5_real); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_io_in_imag = fft_fft_SDFChainRadix22__T_793 ? $signed(fft_fft_SDFChainRadix22__T_799) : $signed(fft_fft_SDFChainRadix22_outputWires_5_imag); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_io_cntr = {{2'd0}, fft_fft_SDFChainRadix22__T_209}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_6_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_7_io_in_real = fft_fft_SDFChainRadix22__T_2110[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_io_in_imag = fft_fft_SDFChainRadix22__T_2114[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_io_cntr = {{1'd0}, fft_fft_SDFChainRadix22__T_216}; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_7_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_clock = fft_fft_SDFChainRadix22_clock;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_reset = fft_fft_SDFChainRadix22_reset;
  assign fft_fft_SDFChainRadix22_sdf_stages_8_io_in_real = fft_fft_SDFChainRadix22__T_2124 ? $signed(fft_fft_SDFChainRadix22_outputWires_7_imag) : $signed(fft_fft_SDFChainRadix22_outputWires_7_real); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_io_in_imag = fft_fft_SDFChainRadix22__T_2124 ? $signed(fft_fft_SDFChainRadix22__T_2130) : $signed(fft_fft_SDFChainRadix22_outputWires_7_imag); // @[SDFChainRadix22.scala 340:23]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_io_cntr = fft_fft_SDFChainRadix22_cntr_wires_0 - fft_fft_SDFChainRadix22__T_220; // @[SDFChainRadix22.scala 224:16]
  assign fft_fft_SDFChainRadix22_sdf_stages_8_io_en = fft_fft_SDFChainRadix22__T_46 | fft_fft_SDFChainRadix22__T_122; // @[SDFChainRadix22.scala 223:14]
  assign fft_fft__T_152 = $signed(fft_fft_io_in_bits_real) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  assign fft_fft__T_153 = $signed(fft_fft_io_in_bits_imag) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  assign fft_fft_io_in_ready = fft_fft_SDFChainRadix22_io_in_ready; // @[SDFFFT.scala 305:23 SDFFFT.scala 309:21]
  assign fft_fft_io_out_valid = fft_fft_SDFChainRadix22_io_out_valid; // @[SDFFFT.scala 306:18 SDFFFT.scala 313:24]
  assign fft_fft_io_out_bits_real = fft_fft_SDFChainRadix22_io_out_bits_real; // @[SDFFFT.scala 306:18 SDFFFT.scala 311:23]
  assign fft_fft_io_out_bits_imag = fft_fft_SDFChainRadix22_io_out_bits_imag; // @[SDFFFT.scala 306:18 SDFFFT.scala 311:23]
  assign fft_fft_io_lastOut = fft_fft_SDFChainRadix22_io_lastOut; // @[SDFFFT.scala 317:20]
  assign fft_fft_io_busy = fft_fft_SDFChainRadix22_io_busy; // @[SDFFFT.scala 320:15]
  assign fft_fft_SDFChainRadix22_clock = fft_fft_clock;
  assign fft_fft_SDFChainRadix22_reset = fft_fft_reset;
  assign fft_fft_SDFChainRadix22_io_in_valid = fft_fft_io_in_valid; // @[SDFFFT.scala 304:27 SDFFFT.scala 309:21]
  assign fft_fft__GEN_526 = fft_fft__T_152[31:14]; // @[SDFFFT.scala 301:31 SDFFFT.scala 309:21]
  assign fft_fft_SDFChainRadix22_io_in_bits_real = fft_fft__GEN_526[15:0]; // @[SDFFFT.scala 301:31 SDFFFT.scala 309:21]
  assign fft_fft__GEN_528 = fft_fft__T_153[31:14]; // @[SDFFFT.scala 302:31 SDFFFT.scala 309:21]
  assign fft_fft_SDFChainRadix22_io_in_bits_imag = fft_fft__GEN_528[15:0]; // @[SDFFFT.scala 302:31 SDFFFT.scala 309:21]
  assign fft_fft_SDFChainRadix22_io_out_ready = fft_fft_io_out_ready; // @[SDFFFT.scala 306:18 SDFFFT.scala 314:28]
  assign fft_fft_SDFChainRadix22_io_lastIn = fft_fft_io_lastIn; // @[SDFFFT.scala 316:23]
  assign fft_Queue__T_read__T_18_addr = fft_Queue_value_1;
  assign fft_Queue__T_read__T_18_data = fft_Queue__T_read[fft_Queue__T_read__T_18_addr]; // @[Decoupled.scala 209:24]
  assign fft_Queue__T_read__T_10_data = fft_Queue_io_enq_bits_read;
  assign fft_Queue__T_read__T_10_addr = fft_Queue_value;
  assign fft_Queue__T_read__T_10_mask = 1'h1;
  assign fft_Queue__T_read__T_10_en = fft_Queue_io_enq_ready & fft_Queue_io_enq_valid;
  assign fft_Queue__T_data__T_18_addr = fft_Queue_value_1;
  assign fft_Queue__T_data__T_18_data = fft_Queue__T_data[fft_Queue__T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign fft_Queue__T_data__T_10_data = fft_Queue_io_enq_bits_data;
  assign fft_Queue__T_data__T_10_addr = fft_Queue_value;
  assign fft_Queue__T_data__T_10_mask = 1'h1;
  assign fft_Queue__T_data__T_10_en = fft_Queue_io_enq_ready & fft_Queue_io_enq_valid;
  assign fft_Queue__T_extra__T_18_addr = fft_Queue_value_1;
  assign fft_Queue__T_extra__T_18_data = fft_Queue__T_extra[fft_Queue__T_extra__T_18_addr]; // @[Decoupled.scala 209:24]
  assign fft_Queue__T_extra__T_10_data = fft_Queue_io_enq_bits_extra;
  assign fft_Queue__T_extra__T_10_addr = fft_Queue_value;
  assign fft_Queue__T_extra__T_10_mask = 1'h1;
  assign fft_Queue__T_extra__T_10_en = fft_Queue_io_enq_ready & fft_Queue_io_enq_valid;
  assign fft_Queue__T_2 = fft_Queue_value == fft_Queue_value_1; // @[Decoupled.scala 214:41]
  assign fft_Queue__T_3 = ~fft_Queue__T_1; // @[Decoupled.scala 215:36]
  assign fft_Queue__T_4 = fft_Queue__T_2 & fft_Queue__T_3; // @[Decoupled.scala 215:33]
  assign fft_Queue__T_5 = fft_Queue__T_2 & fft_Queue__T_1; // @[Decoupled.scala 216:32]
  assign fft_Queue__T_6 = fft_Queue_io_enq_ready & fft_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign fft_Queue__T_8 = fft_Queue_io_deq_ready & fft_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign fft_Queue__T_12 = fft_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign fft_Queue__T_14 = fft_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign fft_Queue__T_15 = fft_Queue__T_6 != fft_Queue__T_8; // @[Decoupled.scala 227:16]
  assign fft_Queue_io_enq_ready = ~fft_Queue__T_5; // @[Decoupled.scala 232:16]
  assign fft_Queue_io_deq_valid = ~fft_Queue__T_4; // @[Decoupled.scala 231:16]
  assign fft_Queue_io_deq_bits_read = fft_Queue__T_read__T_18_data; // @[Decoupled.scala 233:15]
  assign fft_Queue_io_deq_bits_data = fft_Queue__T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign fft_Queue_io_deq_bits_extra = fft_Queue__T_extra__T_18_data; // @[Decoupled.scala 233:15]
  assign fft__T_2 = fft_auto_mem_in_aw_valid & fft_auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign fft__T_4 = ~fft_auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign fft__T_47_ready = fft_Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign fft__T_11 = fft_auto_mem_in_ar_valid ? fft_auto_mem_in_ar_bits_addr : fft_auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign fft__T_45 = fft__T_11[29:2]; // @[RegisterRouter.scala 52:27]
  assign fft__T_1_bits_index = fft__T_45[5:0]; // @[RegisterRouter.scala 37:18 RegisterRouter.scala 52:19]
  assign fft__T_53 = fft__T_1_bits_index == 6'h0; // @[RegisterRouter.scala 59:16]
  assign fft__T_5 = fft__T_47_ready & fft__T_4; // @[RegisterRouter.scala 42:26]
  assign fft__T_171 = fft__T_53 & fft_busy; // @[RegisterRouter.scala 59:16]
  assign fft__T_172_bits_read = fft_Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign fft__T_172_valid = fft_Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign fft__T_175 = ~fft__T_172_bits_read; // @[RegisterRouter.scala 65:29]
  assign fft_auto_mem_in_aw_ready = fft__T_5 & fft_auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign fft_auto_mem_in_w_ready = fft__T_5 & fft_auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign fft_auto_mem_in_b_valid = fft__T_172_valid & fft__T_175; // @[LazyModule.scala 173:31]
  assign fft_auto_mem_in_b_bits_id = fft_Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign fft_auto_mem_in_ar_ready = fft_Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign fft_auto_mem_in_r_valid = fft__T_172_valid & fft__T_172_bits_read; // @[LazyModule.scala 173:31]
  assign fft_auto_mem_in_r_bits_id = fft_Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign fft_auto_mem_in_r_bits_data = fft_Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign fft_auto_stream_in_ready = fft_fft_io_in_ready; // @[LazyModule.scala 173:31]
  assign fft_auto_stream_out_valid = fft_fft_io_out_valid; // @[LazyModule.scala 173:49]
  assign fft_auto_stream_out_bits_data = {fft_fft_io_out_bits_real,fft_fft_io_out_bits_imag}; // @[LazyModule.scala 173:49]
  assign fft_auto_stream_out_bits_last = fft_fft_io_lastOut; // @[LazyModule.scala 173:49]
  assign fft_fft_clock = fft_clock;
  assign fft_fft_reset = fft_reset;
  assign fft_fft_io_in_valid = fft_auto_stream_in_valid; // @[FFTBlock.scala 124:24]
  assign fft_fft_io_in_bits_real = fft_auto_stream_in_bits_data[31:16]; // @[FFTBlock.scala 130:26]
  assign fft_fft_io_in_bits_imag = fft_auto_stream_in_bits_data[15:0]; // @[FFTBlock.scala 129:26]
  assign fft_fft_io_out_ready = fft_auto_stream_out_ready; // @[FFTBlock.scala 137:22]
  assign fft_fft_io_lastIn = fft_auto_stream_in_bits_last; // @[FFTBlock.scala 133:24]
  assign fft_Queue_clock = fft_clock;
  assign fft_Queue_reset = fft_reset;
  assign fft_Queue_io_enq_valid = fft_auto_mem_in_ar_valid | fft__T_2; // @[Decoupled.scala 288:22]
  assign fft_Queue_io_enq_bits_read = fft_auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign fft_Queue_io_enq_bits_data = {{31'd0}, fft__T_171}; // @[Decoupled.scala 289:21]
  assign fft_Queue_io_enq_bits_extra = fft_auto_mem_in_ar_valid ? fft_auto_mem_in_ar_bits_id : fft_auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign fft_Queue_io_deq_ready = fft__T_172_bits_read ? fft_auto_mem_in_r_ready : fft_auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
  assign mag_logMagMux_magModule_Queue__T__T_18_addr = mag_logMagMux_magModule_Queue_value_1;
  assign mag_logMagMux_magModule_Queue__T__T_18_data = mag_logMagMux_magModule_Queue__T[mag_logMagMux_magModule_Queue__T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign mag_logMagMux_magModule_Queue__T__T_10_data = mag_logMagMux_magModule_Queue_io_enq_bits;
  assign mag_logMagMux_magModule_Queue__T__T_10_addr = mag_logMagMux_magModule_Queue_value;
  assign mag_logMagMux_magModule_Queue__T__T_10_mask = 1'h1;
  assign mag_logMagMux_magModule_Queue__T__T_10_en = mag_logMagMux_magModule_Queue_io_enq_ready & mag_logMagMux_magModule_Queue_io_enq_valid;
  assign mag_logMagMux_magModule_Queue__T_2 = mag_logMagMux_magModule_Queue_value == mag_logMagMux_magModule_Queue_value_1; // @[Decoupled.scala 214:41]
  assign mag_logMagMux_magModule_Queue__T_3 = ~mag_logMagMux_magModule_Queue__T_1; // @[Decoupled.scala 215:36]
  assign mag_logMagMux_magModule_Queue__T_4 = mag_logMagMux_magModule_Queue__T_2 & mag_logMagMux_magModule_Queue__T_3; // @[Decoupled.scala 215:33]
  assign mag_logMagMux_magModule_Queue__T_5 = mag_logMagMux_magModule_Queue__T_2 & mag_logMagMux_magModule_Queue__T_1; // @[Decoupled.scala 216:32]
  assign mag_logMagMux_magModule_Queue__T_6 = mag_logMagMux_magModule_Queue_io_enq_ready & mag_logMagMux_magModule_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule_Queue__T_8 = mag_logMagMux_magModule_Queue_io_deq_ready & mag_logMagMux_magModule_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule_Queue__T_12 = mag_logMagMux_magModule_Queue_value + 2'h1; // @[Counter.scala 39:22]
  assign mag_logMagMux_magModule_Queue__T_14 = mag_logMagMux_magModule_Queue_value_1 + 2'h1; // @[Counter.scala 39:22]
  assign mag_logMagMux_magModule_Queue__T_15 = mag_logMagMux_magModule_Queue__T_6 != mag_logMagMux_magModule_Queue__T_8; // @[Decoupled.scala 227:16]
  assign mag_logMagMux_magModule_Queue_io_enq_ready = ~mag_logMagMux_magModule_Queue__T_5; // @[Decoupled.scala 232:16]
  assign mag_logMagMux_magModule_Queue_io_deq_valid = ~mag_logMagMux_magModule_Queue__T_4; // @[Decoupled.scala 231:16]
  assign mag_logMagMux_magModule_Queue_io_deq_bits = mag_logMagMux_magModule_Queue__T__T_18_data; // @[Decoupled.scala 233:15]
  assign mag_logMagMux_magModule_Queue_1__T__T_18_addr = mag_logMagMux_magModule_Queue_1_value_1;
  assign mag_logMagMux_magModule_Queue_1__T__T_18_data = mag_logMagMux_magModule_Queue_1__T[mag_logMagMux_magModule_Queue_1__T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign mag_logMagMux_magModule_Queue_1__T__T_10_data = mag_logMagMux_magModule_Queue_1_io_enq_bits;
  assign mag_logMagMux_magModule_Queue_1__T__T_10_addr = mag_logMagMux_magModule_Queue_1_value;
  assign mag_logMagMux_magModule_Queue_1__T__T_10_mask = 1'h1;
  assign mag_logMagMux_magModule_Queue_1__T__T_10_en = mag_logMagMux_magModule_Queue_1_io_enq_ready & mag_logMagMux_magModule_Queue_1_io_enq_valid;
  assign mag_logMagMux_magModule_Queue_1__T_2 = mag_logMagMux_magModule_Queue_1_value == mag_logMagMux_magModule_Queue_1_value_1; // @[Decoupled.scala 214:41]
  assign mag_logMagMux_magModule_Queue_1__T_3 = ~mag_logMagMux_magModule_Queue_1__T_1; // @[Decoupled.scala 215:36]
  assign mag_logMagMux_magModule_Queue_1__T_4 = mag_logMagMux_magModule_Queue_1__T_2 & mag_logMagMux_magModule_Queue_1__T_3; // @[Decoupled.scala 215:33]
  assign mag_logMagMux_magModule_Queue_1__T_5 = mag_logMagMux_magModule_Queue_1__T_2 & mag_logMagMux_magModule_Queue_1__T_1; // @[Decoupled.scala 216:32]
  assign mag_logMagMux_magModule_Queue_1__T_6 = mag_logMagMux_magModule_Queue_1_io_enq_ready & mag_logMagMux_magModule_Queue_1_io_enq_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule_Queue_1__T_8 = mag_logMagMux_magModule_Queue_1_io_deq_ready & mag_logMagMux_magModule_Queue_1_io_deq_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule_Queue_1__T_12 = mag_logMagMux_magModule_Queue_1_value + 2'h1; // @[Counter.scala 39:22]
  assign mag_logMagMux_magModule_Queue_1__T_14 = mag_logMagMux_magModule_Queue_1_value_1 + 2'h1; // @[Counter.scala 39:22]
  assign mag_logMagMux_magModule_Queue_1__T_15 = mag_logMagMux_magModule_Queue_1__T_6 != mag_logMagMux_magModule_Queue_1__T_8; // @[Decoupled.scala 227:16]
  assign mag_logMagMux_magModule_Queue_1_io_enq_ready = ~mag_logMagMux_magModule_Queue_1__T_5; // @[Decoupled.scala 232:16]
  assign mag_logMagMux_magModule_Queue_1_io_deq_valid = ~mag_logMagMux_magModule_Queue_1__T_4; // @[Decoupled.scala 231:16]
  assign mag_logMagMux_magModule_Queue_1_io_deq_bits = mag_logMagMux_magModule_Queue_1__T__T_18_data; // @[Decoupled.scala 233:15]
  assign mag_logMagMux_magModule__T_2 = mag_logMagMux_magModule_io_in_bits_real[15]; // @[FixedPointTypeClass.scala 224:24]
  assign mag_logMagMux_magModule__T_5 = 16'sh0 - $signed(mag_logMagMux_magModule_io_in_bits_real); // @[FixedPointTypeClass.scala 30:68]
  assign mag_logMagMux_magModule_absInReal = mag_logMagMux_magModule__T_2 ? $signed(mag_logMagMux_magModule__T_5) : $signed(mag_logMagMux_magModule_io_in_bits_real); // @[FixedPointTypeClass.scala 247:8]
  assign mag_logMagMux_magModule__T_6 = mag_logMagMux_magModule_io_in_bits_imag[15]; // @[FixedPointTypeClass.scala 224:24]
  assign mag_logMagMux_magModule__T_9 = 16'sh0 - $signed(mag_logMagMux_magModule_io_in_bits_imag); // @[FixedPointTypeClass.scala 30:68]
  assign mag_logMagMux_magModule_absInImag = mag_logMagMux_magModule__T_6 ? $signed(mag_logMagMux_magModule__T_9) : $signed(mag_logMagMux_magModule_io_in_bits_imag); // @[FixedPointTypeClass.scala 247:8]
  assign mag_logMagMux_magModule__T_10 = $signed(mag_logMagMux_magModule_absInReal) > $signed(mag_logMagMux_magModule_absInImag); // @[FixedPointTypeClass.scala 55:59]
  assign mag_logMagMux_magModule_u = mag_logMagMux_magModule__T_10 ? $signed(mag_logMagMux_magModule_absInReal) : $signed(mag_logMagMux_magModule_absInImag); // @[Order.scala 56:31]
  assign mag_logMagMux_magModule__T_11 = $signed(mag_logMagMux_magModule_absInReal) < $signed(mag_logMagMux_magModule_absInImag); // @[FixedPointTypeClass.scala 53:59]
  assign mag_logMagMux_magModule_v = mag_logMagMux_magModule__T_11 ? $signed(mag_logMagMux_magModule_absInReal) : $signed(mag_logMagMux_magModule_absInImag); // @[Order.scala 55:31]
  assign mag_logMagMux_magModule__T_12 = mag_logMagMux_magModule_v[15:3]; // @[FixedPointTypeClass.scala 117:50]
  assign mag_logMagMux_magModule__GEN_16 = {{3{mag_logMagMux_magModule__T_12[12]}},mag_logMagMux_magModule__T_12}; // @[FixedPointTypeClass.scala 24:22]
  assign mag_logMagMux_magModule__T_15 = mag_logMagMux_magModule_u[15:3]; // @[FixedPointTypeClass.scala 117:50]
  assign mag_logMagMux_magModule__GEN_17 = {{3{mag_logMagMux_magModule__T_15[12]}},mag_logMagMux_magModule__T_15}; // @[FixedPointTypeClass.scala 33:22]
  assign mag_logMagMux_magModule__GEN_18 = {{2{mag_logMagMux_magModule__T_18[14]}},mag_logMagMux_magModule__T_18}; // @[FixedPointTypeClass.scala 24:22]
  assign mag_logMagMux_magModule__T_22 = mag_logMagMux_magModule__T_21[31:14]; // @[FixedPointTypeClass.scala 153:43]
  assign mag_logMagMux_magModule__T_25 = mag_logMagMux_magModule__T_24[31:14]; // @[FixedPointTypeClass.scala 153:43]
  assign mag_logMagMux_magModule__GEN_19 = {{1{mag_logMagMux_magModule_jplMagOp1[16]}},mag_logMagMux_magModule_jplMagOp1}; // @[FixedPointTypeClass.scala 55:59]
  assign mag_logMagMux_magModule__T_33 = $signed(mag_logMagMux_magModule__GEN_19) > $signed(mag_logMagMux_magModule_jplMagOp2); // @[FixedPointTypeClass.scala 55:59]
  assign mag_logMagMux_magModule_jplMag = mag_logMagMux_magModule__T_33 ? $signed({{1{mag_logMagMux_magModule_jplMagOp1[16]}},mag_logMagMux_magModule_jplMagOp1}) : $signed(mag_logMagMux_magModule_jplMagOp2); // @[Order.scala 56:31]
  assign mag_logMagMux_magModule__T_38 = 2'h0 == mag_logMagMux_magModule__T_35; // @[Mux.scala 68:19]
  assign mag_logMagMux_magModule__T_39 = mag_logMagMux_magModule__T_38 ? $signed(mag_logMagMux_magModule_squared_magnitude) : $signed({{1{mag_logMagMux_magModule_jplMag[17]}},mag_logMagMux_magModule_jplMag}); // @[Mux.scala 68:16]
  assign mag_logMagMux_magModule__T_48 = mag_logMagMux_magModule_queueCounter < 2'h3; // @[Skid.scala 35:31]
  assign mag_logMagMux_magModule__T_49 = mag_logMagMux_magModule_queueCounter == 2'h3; // @[Skid.scala 35:68]
  assign mag_logMagMux_magModule__T_50 = mag_logMagMux_magModule__T_49 & mag_logMagMux_magModule_io_out_ready; // @[Skid.scala 35:89]
  assign mag_logMagMux_magModule_skidInData_ready = mag_logMagMux_magModule__T_48 | mag_logMagMux_magModule__T_50; // @[Skid.scala 35:51]
  assign mag_logMagMux_magModule__T_40 = mag_logMagMux_magModule_skidInData_ready & mag_logMagMux_magModule_io_in_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule__GEN_20 = {{1'd0}, mag_logMagMux_magModule__T_40}; // @[Skid.scala 28:34]
  assign mag_logMagMux_magModule__T_41 = mag_logMagMux_magModule_queueCounter + mag_logMagMux_magModule__GEN_20; // @[Skid.scala 28:34]
  assign mag_logMagMux_magModule__T_42 = mag_logMagMux_magModule_io_out_ready & mag_logMagMux_magModule_io_out_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule__GEN_21 = {{2'd0}, mag_logMagMux_magModule__T_42}; // @[Skid.scala 28:47]
  assign mag_logMagMux_magModule__T_43 = mag_logMagMux_magModule__T_41 - mag_logMagMux_magModule__GEN_21; // @[Skid.scala 28:47]
  assign mag_logMagMux_magModule__T_54 = mag_logMagMux_magModule_io_in_ready & mag_logMagMux_magModule_io_in_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule__T_66 = mag_logMagMux_magModule_queueCounter_1 < 2'h3; // @[Skid.scala 35:31]
  assign mag_logMagMux_magModule__T_67 = mag_logMagMux_magModule_queueCounter_1 == 2'h3; // @[Skid.scala 35:68]
  assign mag_logMagMux_magModule__T_68 = mag_logMagMux_magModule__T_67 & mag_logMagMux_magModule_io_out_ready; // @[Skid.scala 35:89]
  assign mag_logMagMux_magModule__T_69 = mag_logMagMux_magModule__T_66 | mag_logMagMux_magModule__T_68; // @[Skid.scala 35:51]
  assign mag_logMagMux_magModule__T_58 = mag_logMagMux_magModule__T_69 & mag_logMagMux_magModule_io_in_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule__GEN_22 = {{1'd0}, mag_logMagMux_magModule__T_58}; // @[Skid.scala 28:34]
  assign mag_logMagMux_magModule__T_59 = mag_logMagMux_magModule_queueCounter_1 + mag_logMagMux_magModule__GEN_22; // @[Skid.scala 28:34]
  assign mag_logMagMux_magModule__T_53_valid = mag_logMagMux_magModule_Queue_1_io_deq_valid; // @[LogMagMuxTypes.scala 220:27 Skid.scala 37:15]
  assign mag_logMagMux_magModule__T_60 = mag_logMagMux_magModule_io_out_ready & mag_logMagMux_magModule__T_53_valid; // @[Decoupled.scala 40:37]
  assign mag_logMagMux_magModule__GEN_23 = {{2'd0}, mag_logMagMux_magModule__T_60}; // @[Skid.scala 28:47]
  assign mag_logMagMux_magModule__T_61 = mag_logMagMux_magModule__T_59 - mag_logMagMux_magModule__GEN_23; // @[Skid.scala 28:47]
  assign mag_logMagMux_magModule_io_in_ready = mag_logMagMux_magModule__T_48 | mag_logMagMux_magModule__T_50; // @[LogMagMuxTypes.scala 215:15]
  assign mag_logMagMux_magModule_io_out_valid = mag_logMagMux_magModule_Queue_io_deq_valid; // @[Skid.scala 37:15]
  assign mag_logMagMux_magModule_io_out_bits = mag_logMagMux_magModule_Queue_io_deq_bits; // @[Skid.scala 38:14]
  assign mag_logMagMux_magModule_io_lastOut = mag_logMagMux_magModule_Queue_1_io_deq_bits; // @[LogMagMuxTypes.scala 225:20]
  assign mag_logMagMux_magModule_Queue_clock = mag_logMagMux_magModule_clock;
  assign mag_logMagMux_magModule_Queue_reset = mag_logMagMux_magModule_reset;
  assign mag_logMagMux_magModule_Queue_io_enq_valid = mag_logMagMux_magModule__T_47; // @[Skid.scala 30:24]
  assign mag_logMagMux_magModule_Queue_io_enq_bits = mag_logMagMux_magModule__T_39[15:0]; // @[LogMagMuxTypes.scala 216:37]
  assign mag_logMagMux_magModule_Queue_io_deq_ready = mag_logMagMux_magModule_io_out_ready; // @[Skid.scala 36:24]
  assign mag_logMagMux_magModule_Queue_1_clock = mag_logMagMux_magModule_clock;
  assign mag_logMagMux_magModule_Queue_1_reset = mag_logMagMux_magModule_reset;
  assign mag_logMagMux_magModule_Queue_1_io_enq_valid = mag_logMagMux_magModule__T_65; // @[Skid.scala 30:24]
  assign mag_logMagMux_magModule_Queue_1_io_enq_bits = mag_logMagMux_magModule__T_57; // @[LogMagMuxTypes.scala 224:44]
  assign mag_logMagMux_magModule_Queue_1_io_deq_ready = mag_logMagMux_magModule_io_out_ready; // @[Skid.scala 36:24]
  assign mag_logMagMux_io_in_ready = mag_logMagMux_magModule_io_in_ready; // @[LogMagMuxGenerator.scala 64:19]
  assign mag_logMagMux_io_out_valid = mag_logMagMux_magModule_io_out_valid; // @[LogMagMuxGenerator.scala 65:10]
  assign mag_logMagMux_io_out_bits = mag_logMagMux_magModule_io_out_bits; // @[LogMagMuxGenerator.scala 65:10]
  assign mag_logMagMux_io_lastOut = mag_logMagMux_magModule_io_lastOut; // @[LogMagMuxGenerator.scala 73:20]
  assign mag_logMagMux_magModule_clock = mag_logMagMux_clock;
  assign mag_logMagMux_magModule_reset = mag_logMagMux_reset;
  assign mag_logMagMux_magModule_io_in_valid = mag_logMagMux_io_in_valid; // @[LogMagMuxGenerator.scala 64:19]
  assign mag_logMagMux_magModule_io_in_bits_real = mag_logMagMux_io_in_bits_real; // @[LogMagMuxGenerator.scala 64:19]
  assign mag_logMagMux_magModule_io_in_bits_imag = mag_logMagMux_io_in_bits_imag; // @[LogMagMuxGenerator.scala 64:19]
  assign mag_logMagMux_magModule_io_lastIn = mag_logMagMux_io_lastIn; // @[LogMagMuxGenerator.scala 72:29]
  assign mag_logMagMux_magModule_io_out_ready = mag_logMagMux_io_out_ready; // @[LogMagMuxGenerator.scala 65:10]
  assign mag_logMagMux_magModule_io_sel = mag_logMagMux_io_sel; // @[LogMagMuxGenerator.scala 68:26]
  assign mag_Queue__T_read__T_18_addr = mag_Queue_value_1;
  assign mag_Queue__T_read__T_18_data = mag_Queue__T_read[mag_Queue__T_read__T_18_addr]; // @[Decoupled.scala 209:24]
  assign mag_Queue__T_read__T_10_data = mag_Queue_io_enq_bits_read;
  assign mag_Queue__T_read__T_10_addr = mag_Queue_value;
  assign mag_Queue__T_read__T_10_mask = 1'h1;
  assign mag_Queue__T_read__T_10_en = mag_Queue_io_enq_ready & mag_Queue_io_enq_valid;
  assign mag_Queue__T_data__T_18_addr = mag_Queue_value_1;
  assign mag_Queue__T_data__T_18_data = mag_Queue__T_data[mag_Queue__T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign mag_Queue__T_data__T_10_data = mag_Queue_io_enq_bits_data;
  assign mag_Queue__T_data__T_10_addr = mag_Queue_value;
  assign mag_Queue__T_data__T_10_mask = 1'h1;
  assign mag_Queue__T_data__T_10_en = mag_Queue_io_enq_ready & mag_Queue_io_enq_valid;
  assign mag_Queue__T_extra__T_18_addr = mag_Queue_value_1;
  assign mag_Queue__T_extra__T_18_data = mag_Queue__T_extra[mag_Queue__T_extra__T_18_addr]; // @[Decoupled.scala 209:24]
  assign mag_Queue__T_extra__T_10_data = mag_Queue_io_enq_bits_extra;
  assign mag_Queue__T_extra__T_10_addr = mag_Queue_value;
  assign mag_Queue__T_extra__T_10_mask = 1'h1;
  assign mag_Queue__T_extra__T_10_en = mag_Queue_io_enq_ready & mag_Queue_io_enq_valid;
  assign mag_Queue__T_2 = mag_Queue_value == mag_Queue_value_1; // @[Decoupled.scala 214:41]
  assign mag_Queue__T_3 = ~mag_Queue__T_1; // @[Decoupled.scala 215:36]
  assign mag_Queue__T_4 = mag_Queue__T_2 & mag_Queue__T_3; // @[Decoupled.scala 215:33]
  assign mag_Queue__T_5 = mag_Queue__T_2 & mag_Queue__T_1; // @[Decoupled.scala 216:32]
  assign mag_Queue__T_6 = mag_Queue_io_enq_ready & mag_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign mag_Queue__T_8 = mag_Queue_io_deq_ready & mag_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign mag_Queue__T_12 = mag_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign mag_Queue__T_14 = mag_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign mag_Queue__T_15 = mag_Queue__T_6 != mag_Queue__T_8; // @[Decoupled.scala 227:16]
  assign mag_Queue_io_enq_ready = ~mag_Queue__T_5; // @[Decoupled.scala 232:16]
  assign mag_Queue_io_deq_valid = ~mag_Queue__T_4; // @[Decoupled.scala 231:16]
  assign mag_Queue_io_deq_bits_read = mag_Queue__T_read__T_18_data; // @[Decoupled.scala 233:15]
  assign mag_Queue_io_deq_bits_data = mag_Queue__T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign mag_Queue_io_deq_bits_extra = mag_Queue__T_extra__T_18_data; // @[Decoupled.scala 233:15]
  assign mag__T_2 = mag_auto_mem_in_aw_valid & mag_auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign mag__T_3 = mag_auto_mem_in_ar_valid | mag__T_2; // @[RegisterRouter.scala 40:26]
  assign mag__T_4 = ~mag_auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign mag__T_47_ready = mag_Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign mag__T_11 = mag_auto_mem_in_ar_valid ? mag_auto_mem_in_ar_bits_addr : mag_auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign mag__T_45 = mag__T_11[29:2]; // @[RegisterRouter.scala 52:27]
  assign mag__T_1_bits_index = mag__T_45[5:0]; // @[RegisterRouter.scala 37:18 RegisterRouter.scala 52:19]
  assign mag__T_53 = mag__T_1_bits_index == 6'h0; // @[RegisterRouter.scala 59:16]
  assign mag__T_5 = mag__T_47_ready & mag__T_4; // @[RegisterRouter.scala 42:26]
  assign mag__T_13 = mag_auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 64:49]
  assign mag__T_14 = 2'h1 << mag__T_13; // @[OneHot.scala 65:12]
  assign mag__T_16 = mag__T_14 | 2'h1; // @[Misc.scala 200:81]
  assign mag__T_17 = mag_auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign mag__T_18 = mag__T_16[1]; // @[Misc.scala 207:26]
  assign mag__T_19 = mag_auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 208:26]
  assign mag__T_20 = ~mag__T_19; // @[Misc.scala 209:20]
  assign mag__T_22 = mag__T_18 & mag__T_20; // @[Misc.scala 213:38]
  assign mag__T_23 = mag__T_17 | mag__T_22; // @[Misc.scala 213:29]
  assign mag__T_25 = mag__T_18 & mag__T_19; // @[Misc.scala 213:38]
  assign mag__T_26 = mag__T_17 | mag__T_25; // @[Misc.scala 213:29]
  assign mag__T_27 = mag__T_16[0]; // @[Misc.scala 207:26]
  assign mag__T_28 = mag_auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 208:26]
  assign mag__T_29 = ~mag__T_28; // @[Misc.scala 209:20]
  assign mag__T_30 = mag__T_20 & mag__T_29; // @[Misc.scala 212:27]
  assign mag__T_31 = mag__T_27 & mag__T_30; // @[Misc.scala 213:38]
  assign mag__T_32 = mag__T_23 | mag__T_31; // @[Misc.scala 213:29]
  assign mag__T_33 = mag__T_20 & mag__T_28; // @[Misc.scala 212:27]
  assign mag__T_34 = mag__T_27 & mag__T_33; // @[Misc.scala 213:38]
  assign mag__T_35 = mag__T_23 | mag__T_34; // @[Misc.scala 213:29]
  assign mag__T_36 = mag__T_19 & mag__T_29; // @[Misc.scala 212:27]
  assign mag__T_37 = mag__T_27 & mag__T_36; // @[Misc.scala 213:38]
  assign mag__T_38 = mag__T_26 | mag__T_37; // @[Misc.scala 213:29]
  assign mag__T_39 = mag__T_19 & mag__T_28; // @[Misc.scala 212:27]
  assign mag__T_40 = mag__T_27 & mag__T_39; // @[Misc.scala 213:38]
  assign mag__T_41 = mag__T_26 | mag__T_40; // @[Misc.scala 213:29]
  assign mag__T_44 = {mag__T_41,mag__T_38,mag__T_35,mag__T_32}; // @[Cat.scala 29:58]
  assign mag__T_46 = mag_auto_mem_in_ar_valid ? mag__T_44 : mag_auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign mag__T_58 = mag__T_46[0]; // @[Bitwise.scala 26:51]
  assign mag__T_59 = mag__T_46[1]; // @[Bitwise.scala 26:51]
  assign mag__T_60 = mag__T_46[2]; // @[Bitwise.scala 26:51]
  assign mag__T_61 = mag__T_46[3]; // @[Bitwise.scala 26:51]
  assign mag__T_63 = mag__T_58 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign mag__T_65 = mag__T_59 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign mag__T_67 = mag__T_60 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign mag__T_69 = mag__T_61 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign mag__T_72 = {mag__T_69,mag__T_67,mag__T_65,mag__T_63}; // @[Cat.scala 29:58]
  assign mag__T_88 = mag__T_72[0]; // @[RegisterRouter.scala 59:16]
  assign mag__T_117 = mag__T_3 & mag__T_47_ready; // @[RegisterRouter.scala 59:16]
  assign mag__T_129 = mag__T_117 & mag__T_4; // @[RegisterRouter.scala 59:16]
  assign mag__T_132 = mag__T_129 & mag__T_53; // @[RegisterRouter.scala 59:16]
  assign mag__T_98 = mag__T_132 & mag__T_88; // @[RegisterRouter.scala 59:16]
  assign mag__T_100 = mag_auto_mem_in_w_bits_data[0]; // @[RegisterRouter.scala 59:16]
  assign mag__T_171 = mag__T_53 & mag_selReg; // @[RegisterRouter.scala 59:16]
  assign mag__T_172_bits_read = mag_Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign mag__T_172_valid = mag_Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign mag__T_175 = ~mag__T_172_bits_read; // @[RegisterRouter.scala 65:29]
  assign mag_auto_mem_in_aw_ready = mag__T_5 & mag_auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign mag_auto_mem_in_w_ready = mag__T_5 & mag_auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign mag_auto_mem_in_b_valid = mag__T_172_valid & mag__T_175; // @[LazyModule.scala 173:31]
  assign mag_auto_mem_in_b_bits_id = mag_Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign mag_auto_mem_in_ar_ready = mag_Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign mag_auto_mem_in_r_valid = mag__T_172_valid & mag__T_172_bits_read; // @[LazyModule.scala 173:31]
  assign mag_auto_mem_in_r_bits_id = mag_Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign mag_auto_mem_in_r_bits_data = mag_Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign mag_auto_master_out_valid = mag_logMagMux_io_out_valid; // @[LazyModule.scala 173:49]
  assign mag_auto_master_out_bits_data = mag_logMagMux_io_out_bits; // @[LazyModule.scala 173:49]
  assign mag_auto_master_out_bits_last = mag_logMagMux_io_lastOut; // @[LazyModule.scala 173:49]
  assign mag_auto_slave_in_ready = mag_logMagMux_io_in_ready; // @[LazyModule.scala 173:31]
  assign mag_logMagMux_clock = mag_clock;
  assign mag_logMagMux_reset = mag_reset;
  assign mag_logMagMux_io_in_valid = mag_auto_slave_in_valid; // @[LogMagMuxDspBlock.scala 87:30]
  assign mag_logMagMux_io_in_bits_real = mag_auto_slave_in_bits_data[31:16]; // @[LogMagMuxDspBlock.scala 88:30]
  assign mag_logMagMux_io_in_bits_imag = mag_auto_slave_in_bits_data[15:0]; // @[LogMagMuxDspBlock.scala 88:30]
  assign mag_logMagMux_io_lastIn = mag_auto_slave_in_bits_last; // @[LogMagMuxDspBlock.scala 91:31]
  assign mag_logMagMux_io_out_ready = mag_auto_master_out_ready; // @[LogMagMuxDspBlock.scala 96:28]
  assign mag_logMagMux_io_sel = {{1'd0}, mag_selReg}; // @[LogMagMuxDspBlock.scala 81:26]
  assign mag_Queue_clock = mag_clock;
  assign mag_Queue_reset = mag_reset;
  assign mag_Queue_io_enq_valid = mag_auto_mem_in_ar_valid | mag__T_2; // @[Decoupled.scala 288:22]
  assign mag_Queue_io_enq_bits_read = mag_auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign mag_Queue_io_enq_bits_data = {{31'd0}, mag__T_171}; // @[Decoupled.scala 289:21]
  assign mag_Queue_io_enq_bits_extra = mag_auto_mem_in_ar_valid ? mag_auto_mem_in_ar_bits_id : mag_auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign mag_Queue_io_deq_ready = mag__T_172_bits_read ? mag_auto_mem_in_r_ready : mag_auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
  assign cfar_cfar_cfarCore_laggWindow_mem__T_423_addr = cfar_cfar_cfarCore_laggWindow_readIdx;
  assign cfar_cfar_cfarCore_laggWindow_mem__T_423_data = cfar_cfar_cfarCore_laggWindow_mem[cfar_cfar_cfarCore_laggWindow_mem__T_423_addr]; // @[CFARUtils.scala 505:26]
  assign cfar_cfar_cfarCore_laggWindow_mem__T_418_data = cfar_cfar_cfarCore_laggWindow_io_in_bits;
  assign cfar_cfar_cfarCore_laggWindow_mem__T_418_addr = cfar_cfar_cfarCore_laggWindow_writeIdxReg;
  assign cfar_cfar_cfarCore_laggWindow_mem__T_418_mask = 1'h1;
  assign cfar_cfar_cfarCore_laggWindow_mem__T_418_en = cfar_cfar_cfarCore_laggWindow_en & cfar_cfar_cfarCore_laggWindow__T_416;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_14_addr = 1'h0;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_14_data = cfar_cfar_cfarCore_laggWindow_outputQueue__T[cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_14_addr]; // @[Decoupled.scala 209:24]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_data = cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_bits;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_addr = 1'h0;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_mask = 1'h1;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_en = cfar_cfar_cfarCore_laggWindow_outputQueue__T_3 ? cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_7 : cfar_cfar_cfarCore_laggWindow_outputQueue__T_6;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T_3 = ~cfar_cfar_cfarCore_laggWindow_outputQueue__T_1; // @[Decoupled.scala 215:36]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T_6 = cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_ready & cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T_8 = cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_ready & cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_7 = cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_ready ? 1'h0 : cfar_cfar_cfarCore_laggWindow_outputQueue__T_6; // @[Decoupled.scala 240:27]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_10 = cfar_cfar_cfarCore_laggWindow_outputQueue__T_3 ? cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_7 : cfar_cfar_cfarCore_laggWindow_outputQueue__T_6; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_9 = cfar_cfar_cfarCore_laggWindow_outputQueue__T_3 ? 1'h0 : cfar_cfar_cfarCore_laggWindow_outputQueue__T_8; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T_11 = cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_10 != cfar_cfar_cfarCore_laggWindow_outputQueue__GEN_9; // @[Decoupled.scala 227:16]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue__T_12 = ~cfar_cfar_cfarCore_laggWindow_outputQueue__T_3; // @[Decoupled.scala 231:19]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_ready = cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_ready | cfar_cfar_cfarCore_laggWindow_outputQueue__T_3; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_valid = cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_valid | cfar_cfar_cfarCore_laggWindow_outputQueue__T_12; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_bits = cfar_cfar_cfarCore_laggWindow_outputQueue__T_3 ? $signed(cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_bits) : $signed(cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_14_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign cfar_cfar_cfarCore_laggWindow__T = cfar_cfar_cfarCore_laggWindow_io_in_ready & cfar_cfar_cfarCore_laggWindow_io_in_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_laggWindow__T_1 = cfar_cfar_cfarCore_laggWindow_last & cfar_cfar_cfarCore_laggWindow_io_out_ready; // @[CFARUtils.scala 511:45]
  assign cfar_cfar_cfarCore_laggWindow_en = cfar_cfar_cfarCore_laggWindow__T | cfar_cfar_cfarCore_laggWindow__T_1; // @[CFARUtils.scala 511:36]
  assign cfar_cfar_cfarCore_laggWindow__T_3 = cfar_cfar_cfarCore_laggWindow_writeIdxReg + 6'h1; // @[CFARUtils.scala 515:21]
  assign cfar_cfar_cfarCore_laggWindow__GEN_140 = {{1'd0}, cfar_cfar_cfarCore_laggWindow__T_3}; // @[CFARUtils.scala 515:27]
  assign cfar_cfar_cfarCore_laggWindow__T_4 = cfar_cfar_cfarCore_laggWindow__GEN_140 >= cfar_cfar_cfarCore_laggWindow_io_depth; // @[CFARUtils.scala 515:27]
  assign cfar_cfar_cfarCore_laggWindow__GEN_141 = {{1'd0}, cfar_cfar_cfarCore_laggWindow_writeIdxReg}; // @[CFARUtils.scala 516:28]
  assign cfar_cfar_cfarCore_laggWindow__T_6 = cfar_cfar_cfarCore_laggWindow__GEN_141 - cfar_cfar_cfarCore_laggWindow_io_depth; // @[CFARUtils.scala 516:28]
  assign cfar_cfar_cfarCore_laggWindow__T_8 = cfar_cfar_cfarCore_laggWindow__T_6 + 7'h1; // @[CFARUtils.scala 516:39]
  assign cfar_cfar_cfarCore_laggWindow__T_10 = 7'h40 + cfar_cfar_cfarCore_laggWindow__GEN_141; // @[CFARUtils.scala 518:27]
  assign cfar_cfar_cfarCore_laggWindow__T_12 = cfar_cfar_cfarCore_laggWindow__T_10 + 7'h1; // @[CFARUtils.scala 518:41]
  assign cfar_cfar_cfarCore_laggWindow__T_14 = cfar_cfar_cfarCore_laggWindow__T_12 - cfar_cfar_cfarCore_laggWindow_io_depth; // @[CFARUtils.scala 518:47]
  assign cfar_cfar_cfarCore_laggWindow__GEN_0 = cfar_cfar_cfarCore_laggWindow__T_4 ? cfar_cfar_cfarCore_laggWindow__T_8 : cfar_cfar_cfarCore_laggWindow__T_14; // @[CFARUtils.scala 515:40]
  assign cfar_cfar_cfarCore_laggWindow__T_16 = cfar_cfar_cfarCore_laggWindow_io_depth - 7'h1; // @[CFARUtils.scala 528:34]
  assign cfar_cfar_cfarCore_laggWindow__T_17 = cfar_cfar_cfarCore_laggWindow__GEN_141 == cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 528:21]
  assign cfar_cfar_cfarCore_laggWindow__T_19 = cfar_cfar_cfarCore_laggWindow__T_17 & cfar_cfar_cfarCore_laggWindow__T; // @[CFARUtils.scala 528:40]
  assign cfar_cfar_cfarCore_laggWindow__GEN_1 = cfar_cfar_cfarCore_laggWindow__T_19 | cfar_cfar_cfarCore_laggWindow_initialInDone; // @[CFARUtils.scala 528:57]
  assign cfar_cfar_cfarCore_laggWindow_fireLastIn = cfar_cfar_cfarCore_laggWindow_io_lastIn & cfar_cfar_cfarCore_laggWindow__T; // @[CFARUtils.scala 531:30]
  assign cfar_cfar_cfarCore_laggWindow__GEN_2 = cfar_cfar_cfarCore_laggWindow_fireLastIn | cfar_cfar_cfarCore_laggWindow_last; // @[CFARUtils.scala 533:21]
  assign cfar_cfar_cfarCore_laggWindow__T_21 = cfar_cfar_cfarCore_laggWindow_io_out_ready & cfar_cfar_cfarCore_laggWindow_io_out_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_laggWindow__T_22 = cfar_cfar_cfarCore_laggWindow_io_depth <= 7'h40; // @[CFARUtils.scala 330:18]
  assign cfar_cfar_cfarCore_laggWindow__T_24 = cfar_cfar_cfarCore_laggWindow__T_22 | cfar_cfar_cfarCore_laggWindow_reset; // @[CFARUtils.scala 330:11]
  assign cfar_cfar_cfarCore_laggWindow__T_25 = ~cfar_cfar_cfarCore_laggWindow__T_24; // @[CFARUtils.scala 330:11]
  assign cfar_cfar_cfarCore_laggWindow__T_33 = 7'h1 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_37 = 7'h2 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_41 = 7'h3 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_45 = 7'h4 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_49 = 7'h5 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_53 = 7'h6 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_57 = 7'h7 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_61 = 7'h8 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_65 = 7'h9 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_69 = 7'ha <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_73 = 7'hb <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_77 = 7'hc <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_81 = 7'hd <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_85 = 7'he <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_89 = 7'hf <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_93 = 7'h10 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_97 = 7'h11 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_101 = 7'h12 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_105 = 7'h13 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_109 = 7'h14 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_113 = 7'h15 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_117 = 7'h16 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_121 = 7'h17 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_125 = 7'h18 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_129 = 7'h19 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_133 = 7'h1a <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_137 = 7'h1b <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_141 = 7'h1c <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_145 = 7'h1d <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_149 = 7'h1e <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_153 = 7'h1f <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_157 = 7'h20 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_161 = 7'h21 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_165 = 7'h22 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_169 = 7'h23 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_173 = 7'h24 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_177 = 7'h25 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_181 = 7'h26 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_185 = 7'h27 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_189 = 7'h28 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_193 = 7'h29 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_197 = 7'h2a <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_201 = 7'h2b <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_205 = 7'h2c <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_209 = 7'h2d <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_213 = 7'h2e <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_217 = 7'h2f <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_221 = 7'h30 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_225 = 7'h31 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_229 = 7'h32 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_233 = 7'h33 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_237 = 7'h34 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_241 = 7'h35 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_245 = 7'h36 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_249 = 7'h37 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_253 = 7'h38 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_257 = 7'h39 <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_261 = 7'h3a <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_265 = 7'h3b <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_269 = 7'h3c <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_273 = 7'h3d <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_277 = 7'h3e <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_281 = 7'h3f <= cfar_cfar_cfarCore_laggWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_laggWindow__T_284 = cfar_cfar_cfarCore_laggWindow__T_281 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_285 = cfar_cfar_cfarCore_laggWindow__T_277 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_286 = cfar_cfar_cfarCore_laggWindow__T_273 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_287 = cfar_cfar_cfarCore_laggWindow__T_269 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_288 = cfar_cfar_cfarCore_laggWindow__T_265 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_289 = cfar_cfar_cfarCore_laggWindow__T_261 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_290 = cfar_cfar_cfarCore_laggWindow__T_257 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_291 = cfar_cfar_cfarCore_laggWindow__T_253 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_292 = cfar_cfar_cfarCore_laggWindow__T_249 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_293 = cfar_cfar_cfarCore_laggWindow__T_245 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_294 = cfar_cfar_cfarCore_laggWindow__T_241 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_295 = cfar_cfar_cfarCore_laggWindow__T_237 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_296 = cfar_cfar_cfarCore_laggWindow__T_233 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_297 = cfar_cfar_cfarCore_laggWindow__T_229 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_298 = cfar_cfar_cfarCore_laggWindow__T_225 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_299 = cfar_cfar_cfarCore_laggWindow__T_221 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_300 = cfar_cfar_cfarCore_laggWindow__T_217 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_301 = cfar_cfar_cfarCore_laggWindow__T_213 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_302 = cfar_cfar_cfarCore_laggWindow__T_209 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_303 = cfar_cfar_cfarCore_laggWindow__T_205 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_304 = cfar_cfar_cfarCore_laggWindow__T_201 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_305 = cfar_cfar_cfarCore_laggWindow__T_197 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_306 = cfar_cfar_cfarCore_laggWindow__T_193 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_307 = cfar_cfar_cfarCore_laggWindow__T_189 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_308 = cfar_cfar_cfarCore_laggWindow__T_185 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_309 = cfar_cfar_cfarCore_laggWindow__T_181 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_310 = cfar_cfar_cfarCore_laggWindow__T_177 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_311 = cfar_cfar_cfarCore_laggWindow__T_173 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_312 = cfar_cfar_cfarCore_laggWindow__T_169 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_313 = cfar_cfar_cfarCore_laggWindow__T_165 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_314 = cfar_cfar_cfarCore_laggWindow__T_161 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_315 = cfar_cfar_cfarCore_laggWindow__T_157 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_316 = cfar_cfar_cfarCore_laggWindow__T_153 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_317 = cfar_cfar_cfarCore_laggWindow__T_149 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_318 = cfar_cfar_cfarCore_laggWindow__T_145 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_319 = cfar_cfar_cfarCore_laggWindow__T_141 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_320 = cfar_cfar_cfarCore_laggWindow__T_137 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_321 = cfar_cfar_cfarCore_laggWindow__T_133 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_322 = cfar_cfar_cfarCore_laggWindow__T_129 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_323 = cfar_cfar_cfarCore_laggWindow__T_125 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_324 = cfar_cfar_cfarCore_laggWindow__T_121 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_325 = cfar_cfar_cfarCore_laggWindow__T_117 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_326 = cfar_cfar_cfarCore_laggWindow__T_113 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_327 = cfar_cfar_cfarCore_laggWindow__T_109 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_328 = cfar_cfar_cfarCore_laggWindow__T_105 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_329 = cfar_cfar_cfarCore_laggWindow__T_101 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_330 = cfar_cfar_cfarCore_laggWindow__T_97 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_331 = cfar_cfar_cfarCore_laggWindow__T_93 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_332 = cfar_cfar_cfarCore_laggWindow__T_89 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_333 = cfar_cfar_cfarCore_laggWindow__T_85 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_334 = cfar_cfar_cfarCore_laggWindow__T_81 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_335 = cfar_cfar_cfarCore_laggWindow__T_77 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_336 = cfar_cfar_cfarCore_laggWindow__T_73 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_337 = cfar_cfar_cfarCore_laggWindow__T_69 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_338 = cfar_cfar_cfarCore_laggWindow__T_65 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_339 = cfar_cfar_cfarCore_laggWindow__T_61 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_340 = cfar_cfar_cfarCore_laggWindow__T_57 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_341 = cfar_cfar_cfarCore_laggWindow__T_53 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_342 = cfar_cfar_cfarCore_laggWindow__T_49 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_343 = cfar_cfar_cfarCore_laggWindow__T_45 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_344 = cfar_cfar_cfarCore_laggWindow__T_41 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_345 = cfar_cfar_cfarCore_laggWindow__T_37 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_346 = cfar_cfar_cfarCore_laggWindow__T_33 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggWindow__T_414 = cfar_cfar_cfarCore_laggWindow__T_16[5:0];
  assign cfar_cfar_cfarCore_laggWindow__GEN_68 = 6'h1 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_349 : cfar_cfar_cfarCore_laggWindow__T_348; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_69 = 6'h2 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_350 : cfar_cfar_cfarCore_laggWindow__GEN_68; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_70 = 6'h3 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_351 : cfar_cfar_cfarCore_laggWindow__GEN_69; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_71 = 6'h4 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_352 : cfar_cfar_cfarCore_laggWindow__GEN_70; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_72 = 6'h5 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_353 : cfar_cfar_cfarCore_laggWindow__GEN_71; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_73 = 6'h6 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_354 : cfar_cfar_cfarCore_laggWindow__GEN_72; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_74 = 6'h7 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_355 : cfar_cfar_cfarCore_laggWindow__GEN_73; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_75 = 6'h8 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_356 : cfar_cfar_cfarCore_laggWindow__GEN_74; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_76 = 6'h9 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_357 : cfar_cfar_cfarCore_laggWindow__GEN_75; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_77 = 6'ha == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_358 : cfar_cfar_cfarCore_laggWindow__GEN_76; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_78 = 6'hb == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_359 : cfar_cfar_cfarCore_laggWindow__GEN_77; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_79 = 6'hc == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_360 : cfar_cfar_cfarCore_laggWindow__GEN_78; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_80 = 6'hd == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_361 : cfar_cfar_cfarCore_laggWindow__GEN_79; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_81 = 6'he == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_362 : cfar_cfar_cfarCore_laggWindow__GEN_80; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_82 = 6'hf == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_363 : cfar_cfar_cfarCore_laggWindow__GEN_81; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_83 = 6'h10 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_364 : cfar_cfar_cfarCore_laggWindow__GEN_82; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_84 = 6'h11 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_365 : cfar_cfar_cfarCore_laggWindow__GEN_83; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_85 = 6'h12 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_366 : cfar_cfar_cfarCore_laggWindow__GEN_84; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_86 = 6'h13 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_367 : cfar_cfar_cfarCore_laggWindow__GEN_85; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_87 = 6'h14 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_368 : cfar_cfar_cfarCore_laggWindow__GEN_86; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_88 = 6'h15 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_369 : cfar_cfar_cfarCore_laggWindow__GEN_87; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_89 = 6'h16 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_370 : cfar_cfar_cfarCore_laggWindow__GEN_88; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_90 = 6'h17 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_371 : cfar_cfar_cfarCore_laggWindow__GEN_89; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_91 = 6'h18 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_372 : cfar_cfar_cfarCore_laggWindow__GEN_90; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_92 = 6'h19 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_373 : cfar_cfar_cfarCore_laggWindow__GEN_91; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_93 = 6'h1a == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_374 : cfar_cfar_cfarCore_laggWindow__GEN_92; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_94 = 6'h1b == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_375 : cfar_cfar_cfarCore_laggWindow__GEN_93; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_95 = 6'h1c == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_376 : cfar_cfar_cfarCore_laggWindow__GEN_94; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_96 = 6'h1d == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_377 : cfar_cfar_cfarCore_laggWindow__GEN_95; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_97 = 6'h1e == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_378 : cfar_cfar_cfarCore_laggWindow__GEN_96; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_98 = 6'h1f == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_379 : cfar_cfar_cfarCore_laggWindow__GEN_97; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_99 = 6'h20 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_380 : cfar_cfar_cfarCore_laggWindow__GEN_98; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_100 = 6'h21 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_381 : cfar_cfar_cfarCore_laggWindow__GEN_99; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_101 = 6'h22 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_382 : cfar_cfar_cfarCore_laggWindow__GEN_100; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_102 = 6'h23 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_383 : cfar_cfar_cfarCore_laggWindow__GEN_101; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_103 = 6'h24 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_384 : cfar_cfar_cfarCore_laggWindow__GEN_102; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_104 = 6'h25 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_385 : cfar_cfar_cfarCore_laggWindow__GEN_103; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_105 = 6'h26 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_386 : cfar_cfar_cfarCore_laggWindow__GEN_104; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_106 = 6'h27 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_387 : cfar_cfar_cfarCore_laggWindow__GEN_105; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_107 = 6'h28 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_388 : cfar_cfar_cfarCore_laggWindow__GEN_106; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_108 = 6'h29 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_389 : cfar_cfar_cfarCore_laggWindow__GEN_107; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_109 = 6'h2a == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_390 : cfar_cfar_cfarCore_laggWindow__GEN_108; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_110 = 6'h2b == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_391 : cfar_cfar_cfarCore_laggWindow__GEN_109; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_111 = 6'h2c == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_392 : cfar_cfar_cfarCore_laggWindow__GEN_110; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_112 = 6'h2d == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_393 : cfar_cfar_cfarCore_laggWindow__GEN_111; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_113 = 6'h2e == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_394 : cfar_cfar_cfarCore_laggWindow__GEN_112; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_114 = 6'h2f == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_395 : cfar_cfar_cfarCore_laggWindow__GEN_113; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_115 = 6'h30 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_396 : cfar_cfar_cfarCore_laggWindow__GEN_114; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_116 = 6'h31 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_397 : cfar_cfar_cfarCore_laggWindow__GEN_115; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_117 = 6'h32 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_398 : cfar_cfar_cfarCore_laggWindow__GEN_116; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_118 = 6'h33 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_399 : cfar_cfar_cfarCore_laggWindow__GEN_117; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_119 = 6'h34 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_400 : cfar_cfar_cfarCore_laggWindow__GEN_118; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_120 = 6'h35 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_401 : cfar_cfar_cfarCore_laggWindow__GEN_119; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_121 = 6'h36 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_402 : cfar_cfar_cfarCore_laggWindow__GEN_120; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_122 = 6'h37 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_403 : cfar_cfar_cfarCore_laggWindow__GEN_121; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_123 = 6'h38 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_404 : cfar_cfar_cfarCore_laggWindow__GEN_122; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_124 = 6'h39 == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_405 : cfar_cfar_cfarCore_laggWindow__GEN_123; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_125 = 6'h3a == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_406 : cfar_cfar_cfarCore_laggWindow__GEN_124; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_126 = 6'h3b == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_407 : cfar_cfar_cfarCore_laggWindow__GEN_125; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_127 = 6'h3c == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_408 : cfar_cfar_cfarCore_laggWindow__GEN_126; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_128 = 6'h3d == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_409 : cfar_cfar_cfarCore_laggWindow__GEN_127; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_129 = 6'h3e == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_410 : cfar_cfar_cfarCore_laggWindow__GEN_128; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__GEN_130 = 6'h3f == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_411 : cfar_cfar_cfarCore_laggWindow__GEN_129; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow_resetAll = cfar_cfar_cfarCore_laggWindow__GEN_130 & cfar_cfar_cfarCore_laggWindow__T_21; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_laggWindow__T_416 = ~cfar_cfar_cfarCore_laggWindow_resetAll; // @[CFARUtils.scala 544:15]
  assign cfar_cfar_cfarCore_laggWindow__T_417 = cfar_cfar_cfarCore_laggWindow_en & cfar_cfar_cfarCore_laggWindow__T_416; // @[CFARUtils.scala 544:12]
  assign cfar_cfar_cfarCore_laggWindow__T_419 = cfar_cfar_cfarCore_laggWindow_writeIdxReg < 6'h3f; // @[CFARUtils.scala 546:36]
  assign cfar_cfar_cfarCore_laggWindow__T_431 = ~cfar_cfar_cfarCore_laggWindow_initialInDone; // @[CFARUtils.scala 554:42]
  assign cfar_cfar_cfarCore_laggWindow__T_433 = ~cfar_cfar_cfarCore_laggWindow_last; // @[CFARUtils.scala 555:36]
  assign cfar_cfar_cfarCore_laggWindow__T_437 = cfar_cfar_cfarCore_laggWindow_io_out_ready & cfar_cfar_cfarCore_laggWindow__T_433; // @[CFARUtils.scala 559:52]
  assign cfar_cfar_cfarCore_laggWindow__T_439 = cfar_cfar_cfarCore_laggWindow_initialInDone & cfar_cfar_cfarCore_laggWindow_io_in_valid; // @[CFARUtils.scala 568:33]
  assign cfar_cfar_cfarCore_laggWindow__T_440 = cfar_cfar_cfarCore_laggWindow_last & cfar_cfar_cfarCore_laggWindow_en; // @[CFARUtils.scala 568:57]
  assign cfar_cfar_cfarCore_laggWindow_readIdx = cfar_cfar_cfarCore_laggWindow__GEN_0[5:0]; // @[CFARUtils.scala 506:27 CFARUtils.scala 516:13 CFARUtils.scala 518:13]
  assign cfar_cfar_cfarCore_laggWindow_io_in_ready = cfar_cfar_cfarCore_laggWindow__T_431 | cfar_cfar_cfarCore_laggWindow__T_437; // @[CFARUtils.scala 559:18]
  assign cfar_cfar_cfarCore_laggWindow_io_out_valid = cfar_cfar_cfarCore_laggWindow__T_439 | cfar_cfar_cfarCore_laggWindow__T_440; // @[CFARUtils.scala 568:16]
  assign cfar_cfar_cfarCore_laggWindow_io_out_bits = cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_bits; // @[CFARUtils.scala 565:16]
  assign cfar_cfar_cfarCore_laggWindow_io_lastOut = 6'h3f == cfar_cfar_cfarCore_laggWindow__T_414 ? cfar_cfar_cfarCore_laggWindow__T_411 : cfar_cfar_cfarCore_laggWindow__GEN_129; // @[CFARUtils.scala 567:16]
  assign cfar_cfar_cfarCore_laggWindow_io_memFull = cfar_cfar_cfarCore_laggWindow_initialInDone & cfar_cfar_cfarCore_laggWindow__T_433; // @[CFARUtils.scala 555:16]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_clock = cfar_cfar_cfarCore_laggWindow_clock;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_reset = cfar_cfar_cfarCore_laggWindow_reset;
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_valid = cfar_cfar_cfarCore_laggWindow_validPrev; // @[CFARUtils.scala 550:28]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_io_enq_bits = cfar_cfar_cfarCore_laggWindow__T_426; // @[CFARUtils.scala 551:27]
  assign cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_ready = cfar_cfar_cfarCore_laggWindow__T | cfar_cfar_cfarCore_laggWindow__T_1; // @[CFARUtils.scala 552:28]
  assign cfar_cfar_cfarCore_laggGuard__T_1 = cfar_cfar_cfarCore_laggGuard_io_in_ready & cfar_cfar_cfarCore_laggGuard_io_in_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_laggGuard__T_2 = cfar_cfar_cfarCore_laggGuard_last & cfar_cfar_cfarCore_laggGuard_io_out_ready; // @[CFARUtils.scala 385:34]
  assign cfar_cfar_cfarCore_laggGuard_en = cfar_cfar_cfarCore_laggGuard__T_1 | cfar_cfar_cfarCore_laggGuard__T_2; // @[CFARUtils.scala 385:25]
  assign cfar_cfar_cfarCore_laggGuard__T_3 = cfar_cfar_cfarCore_laggGuard_io_depth <= 4'h8; // @[CFARUtils.scala 345:18]
  assign cfar_cfar_cfarCore_laggGuard__T_5 = cfar_cfar_cfarCore_laggGuard__T_3 | cfar_cfar_cfarCore_laggGuard_reset; // @[CFARUtils.scala 345:11]
  assign cfar_cfar_cfarCore_laggGuard__T_6 = ~cfar_cfar_cfarCore_laggGuard__T_5; // @[CFARUtils.scala 345:11]
  assign cfar_cfar_cfarCore_laggGuard__T_8 = cfar_cfar_cfarCore_laggGuard_io_depth - 4'h1; // @[CFARUtils.scala 350:87]
  assign cfar_cfar_cfarCore_laggGuard__T_9 = 1'h1; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_13 = 4'h1 <= cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_14 = cfar_cfar_cfarCore_laggGuard__T_13; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_laggGuard__T_17 = 4'h2 <= cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_18 = cfar_cfar_cfarCore_laggGuard__T_17; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_laggGuard__T_21 = 4'h3 <= cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_22 = cfar_cfar_cfarCore_laggGuard__T_21; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_laggGuard__T_25 = 4'h4 <= cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_26 = cfar_cfar_cfarCore_laggGuard__T_25; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_laggGuard__T_29 = 4'h5 <= cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_30 = cfar_cfar_cfarCore_laggGuard__T_29; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_laggGuard__T_33 = 4'h6 <= cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_34 = cfar_cfar_cfarCore_laggGuard__T_33; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_laggGuard__T_37 = 4'h7 <= cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_laggGuard__T_38 = cfar_cfar_cfarCore_laggGuard__T_37; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_laggGuard__T_39 = cfar_cfar_cfarCore_laggGuard__T_38 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_40 = cfar_cfar_cfarCore_laggGuard__T_34 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_41 = cfar_cfar_cfarCore_laggGuard__T_30 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_42 = cfar_cfar_cfarCore_laggGuard__T_26 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_43 = cfar_cfar_cfarCore_laggGuard__T_22 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_44 = cfar_cfar_cfarCore_laggGuard__T_18 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_45 = cfar_cfar_cfarCore_laggGuard__T_14 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_46 = cfar_cfar_cfarCore_laggGuard__T_9 & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_57 = cfar_cfar_cfarCore_laggGuard__T_8[2:0];
  assign cfar_cfar_cfarCore_laggGuard__T_59 = cfar_cfar_cfarCore_laggGuard_io_lastIn & cfar_cfar_cfarCore_laggGuard__T_1; // @[CFARUtils.scala 392:19]
  assign cfar_cfar_cfarCore_laggGuard__GEN_8 = cfar_cfar_cfarCore_laggGuard__T_59 | cfar_cfar_cfarCore_laggGuard_last; // @[CFARUtils.scala 392:36]
  assign cfar_cfar_cfarCore_laggGuard__T_62 = cfar_cfar_cfarCore_laggGuard_cntIn + 4'h1; // @[CFARUtils.scala 397:20]
  assign cfar_cfar_cfarCore_laggGuard__T_63 = cfar_cfar_cfarCore_laggGuard_io_depth > 4'h1; // @[CFARUtils.scala 400:18]
  assign cfar_cfar_cfarCore_laggGuard__T_66 = cfar_cfar_cfarCore_laggGuard_cntIn == cfar_cfar_cfarCore_laggGuard__T_8; // @[CFARUtils.scala 401:17]
  assign cfar_cfar_cfarCore_laggGuard__T_68 = cfar_cfar_cfarCore_laggGuard__T_66 & cfar_cfar_cfarCore_laggGuard__T_1; // @[CFARUtils.scala 401:36]
  assign cfar_cfar_cfarCore_laggGuard__GEN_10 = cfar_cfar_cfarCore_laggGuard__T_68 | cfar_cfar_cfarCore_laggGuard_InitialInDone; // @[CFARUtils.scala 401:53]
  assign cfar_cfar_cfarCore_laggGuard__T_70 = cfar_cfar_cfarCore_laggGuard_io_depth == 4'h1; // @[CFARUtils.scala 406:36]
  assign cfar_cfar_cfarCore_laggGuard__T_71 = cfar_cfar_cfarCore_laggGuard__T_1 & cfar_cfar_cfarCore_laggGuard__T_70; // @[CFARUtils.scala 406:24]
  assign cfar_cfar_cfarCore_laggGuard__GEN_11 = cfar_cfar_cfarCore_laggGuard__T_71 | cfar_cfar_cfarCore_laggGuard_InitialInDone; // @[CFARUtils.scala 406:45]
  assign cfar_cfar_cfarCore_laggGuard__T_73 = cfar_cfar_cfarCore_laggGuard_io_out_ready & cfar_cfar_cfarCore_laggGuard_io_out_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_laggGuard__T_112 = cfar_cfar_cfarCore_laggGuard__T_37 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_113 = cfar_cfar_cfarCore_laggGuard__T_33 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_114 = cfar_cfar_cfarCore_laggGuard__T_29 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_115 = cfar_cfar_cfarCore_laggGuard__T_25 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_116 = cfar_cfar_cfarCore_laggGuard__T_21 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_117 = cfar_cfar_cfarCore_laggGuard__T_17 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__T_118 = cfar_cfar_cfarCore_laggGuard__T_13 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_laggGuard__GEN_22 = 3'h1 == cfar_cfar_cfarCore_laggGuard__T_57 ? cfar_cfar_cfarCore_laggGuard__T_121 : cfar_cfar_cfarCore_laggGuard__T_120; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__GEN_23 = 3'h2 == cfar_cfar_cfarCore_laggGuard__T_57 ? cfar_cfar_cfarCore_laggGuard__T_122 : cfar_cfar_cfarCore_laggGuard__GEN_22; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__GEN_24 = 3'h3 == cfar_cfar_cfarCore_laggGuard__T_57 ? cfar_cfar_cfarCore_laggGuard__T_123 : cfar_cfar_cfarCore_laggGuard__GEN_23; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__GEN_25 = 3'h4 == cfar_cfar_cfarCore_laggGuard__T_57 ? cfar_cfar_cfarCore_laggGuard__T_124 : cfar_cfar_cfarCore_laggGuard__GEN_24; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__GEN_26 = 3'h5 == cfar_cfar_cfarCore_laggGuard__T_57 ? cfar_cfar_cfarCore_laggGuard__T_125 : cfar_cfar_cfarCore_laggGuard__GEN_25; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__GEN_27 = 3'h6 == cfar_cfar_cfarCore_laggGuard__T_57 ? cfar_cfar_cfarCore_laggGuard__T_126 : cfar_cfar_cfarCore_laggGuard__GEN_26; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__GEN_28 = 3'h7 == cfar_cfar_cfarCore_laggGuard__T_57 ? cfar_cfar_cfarCore_laggGuard__T_127 : cfar_cfar_cfarCore_laggGuard__GEN_27; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__T_132 = cfar_cfar_cfarCore_laggGuard__GEN_28 & cfar_cfar_cfarCore_laggGuard__T_73; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_laggGuard__T_134 = ~cfar_cfar_cfarCore_laggGuard_InitialInDone; // @[CFARUtils.scala 420:36]
  assign cfar_cfar_cfarCore_laggGuard__T_136 = ~cfar_cfar_cfarCore_laggGuard_last; // @[CFARUtils.scala 421:36]
  assign cfar_cfar_cfarCore_laggGuard__T_138 = cfar_cfar_cfarCore_laggGuard_io_depth == 4'h0; // @[CFARUtils.scala 426:37]
  assign cfar_cfar_cfarCore_laggGuard__T_141 = cfar_cfar_cfarCore_laggGuard_io_out_ready & cfar_cfar_cfarCore_laggGuard__T_136; // @[CFARUtils.scala 426:91]
  assign cfar_cfar_cfarCore_laggGuard__T_142 = cfar_cfar_cfarCore_laggGuard__T_134 | cfar_cfar_cfarCore_laggGuard__T_141; // @[CFARUtils.scala 426:75]
  assign cfar_cfar_cfarCore_laggGuard__GEN_33 = 3'h1 == cfar_cfar_cfarCore_laggGuard__T_57 ? $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_1) : $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_0); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_laggGuard__GEN_34 = 3'h2 == cfar_cfar_cfarCore_laggGuard__T_57 ? $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_2) : $signed(cfar_cfar_cfarCore_laggGuard__GEN_33); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_laggGuard__GEN_35 = 3'h3 == cfar_cfar_cfarCore_laggGuard__T_57 ? $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_3) : $signed(cfar_cfar_cfarCore_laggGuard__GEN_34); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_laggGuard__GEN_36 = 3'h4 == cfar_cfar_cfarCore_laggGuard__T_57 ? $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_4) : $signed(cfar_cfar_cfarCore_laggGuard__GEN_35); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_laggGuard__GEN_37 = 3'h5 == cfar_cfar_cfarCore_laggGuard__T_57 ? $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_5) : $signed(cfar_cfar_cfarCore_laggGuard__GEN_36); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_laggGuard__GEN_38 = 3'h6 == cfar_cfar_cfarCore_laggGuard__T_57 ? $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_6) : $signed(cfar_cfar_cfarCore_laggGuard__GEN_37); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_laggGuard__GEN_39 = 3'h7 == cfar_cfar_cfarCore_laggGuard__T_57 ? $signed(cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_7) : $signed(cfar_cfar_cfarCore_laggGuard__GEN_38); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_laggGuard__T_151 = cfar_cfar_cfarCore_laggGuard_InitialInDone & cfar_cfar_cfarCore_laggGuard_io_in_valid; // @[CFARUtils.scala 436:70]
  assign cfar_cfar_cfarCore_laggGuard__T_152 = cfar_cfar_cfarCore_laggGuard_last & cfar_cfar_cfarCore_laggGuard_en; // @[CFARUtils.scala 436:94]
  assign cfar_cfar_cfarCore_laggGuard__T_153 = cfar_cfar_cfarCore_laggGuard__T_151 | cfar_cfar_cfarCore_laggGuard__T_152; // @[CFARUtils.scala 436:85]
  assign cfar_cfar_cfarCore_laggGuard_io_in_ready = cfar_cfar_cfarCore_laggGuard__T_138 ? cfar_cfar_cfarCore_laggGuard_io_out_ready : cfar_cfar_cfarCore_laggGuard__T_142; // @[CFARUtils.scala 426:20]
  assign cfar_cfar_cfarCore_laggGuard_io_out_valid = cfar_cfar_cfarCore_laggGuard__T_138 ? cfar_cfar_cfarCore_laggGuard_io_in_valid : cfar_cfar_cfarCore_laggGuard__T_153; // @[CFARUtils.scala 436:18]
  assign cfar_cfar_cfarCore_laggGuard_io_out_bits = cfar_cfar_cfarCore_laggGuard__T_138 ? $signed(cfar_cfar_cfarCore_laggGuard_io_in_bits) : $signed(cfar_cfar_cfarCore_laggGuard__GEN_39); // @[CFARUtils.scala 433:18]
  assign cfar_cfar_cfarCore_laggGuard_io_lastOut = cfar_cfar_cfarCore_laggGuard__T_138 ? cfar_cfar_cfarCore_laggGuard__T_59 : cfar_cfar_cfarCore_laggGuard__GEN_28; // @[CFARUtils.scala 435:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_0 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_0; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_1 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_1; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_2 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_2; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_3 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_3; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_4 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_4; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_5 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_5; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_6 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_6; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_laggGuard_io_parallelOut_7 = cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_7; // @[CFARUtils.scala 434:18]
  assign cfar_cfar_cfarCore_cellUnderTest__T_1 = cfar_cfar_cfarCore_cellUnderTest_io_in_ready & cfar_cfar_cfarCore_cellUnderTest_io_in_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_cellUnderTest__T_2 = ~cfar_cfar_cfarCore_cellUnderTest_initialInDone; // @[CFARUtils.scala 457:25]
  assign cfar_cfar_cfarCore_cellUnderTest__T_3 = cfar_cfar_cfarCore_cellUnderTest__T_1 & cfar_cfar_cfarCore_cellUnderTest__T_2; // @[CFARUtils.scala 457:22]
  assign cfar_cfar_cfarCore_cellUnderTest__GEN_0 = cfar_cfar_cfarCore_cellUnderTest__T_3 | cfar_cfar_cfarCore_cellUnderTest_initialInDone; // @[CFARUtils.scala 457:41]
  assign cfar_cfar_cfarCore_cellUnderTest__T_5 = cfar_cfar_cfarCore_cellUnderTest_last & cfar_cfar_cfarCore_cellUnderTest_io_out_ready; // @[CFARUtils.scala 461:34]
  assign cfar_cfar_cfarCore_cellUnderTest_en = cfar_cfar_cfarCore_cellUnderTest__T_1 | cfar_cfar_cfarCore_cellUnderTest__T_5; // @[CFARUtils.scala 461:25]
  assign cfar_cfar_cfarCore_cellUnderTest__T_7 = cfar_cfar_cfarCore_cellUnderTest_io_lastIn & cfar_cfar_cfarCore_cellUnderTest__T_1; // @[CFARUtils.scala 468:19]
  assign cfar_cfar_cfarCore_cellUnderTest__GEN_2 = cfar_cfar_cfarCore_cellUnderTest__T_7 | cfar_cfar_cfarCore_cellUnderTest_last; // @[CFARUtils.scala 468:36]
  assign cfar_cfar_cfarCore_cellUnderTest__T_9 = cfar_cfar_cfarCore_cellUnderTest_lastOut & cfar_cfar_cfarCore_cellUnderTest_io_out_ready; // @[CFARUtils.scala 475:17]
  assign cfar_cfar_cfarCore_cellUnderTest__T_11 = ~cfar_cfar_cfarCore_cellUnderTest_last; // @[CFARUtils.scala 480:55]
  assign cfar_cfar_cfarCore_cellUnderTest__T_12 = cfar_cfar_cfarCore_cellUnderTest_io_out_ready & cfar_cfar_cfarCore_cellUnderTest__T_11; // @[CFARUtils.scala 480:52]
  assign cfar_cfar_cfarCore_cellUnderTest__T_14 = cfar_cfar_cfarCore_cellUnderTest_initialInDone & cfar_cfar_cfarCore_cellUnderTest_io_in_valid; // @[CFARUtils.scala 483:35]
  assign cfar_cfar_cfarCore_cellUnderTest__T_15 = cfar_cfar_cfarCore_cellUnderTest_last & cfar_cfar_cfarCore_cellUnderTest_en; // @[CFARUtils.scala 483:59]
  assign cfar_cfar_cfarCore_cellUnderTest_io_in_ready = cfar_cfar_cfarCore_cellUnderTest__T_2 | cfar_cfar_cfarCore_cellUnderTest__T_12; // @[CFARUtils.scala 480:18]
  assign cfar_cfar_cfarCore_cellUnderTest_io_out_valid = cfar_cfar_cfarCore_cellUnderTest__T_14 | cfar_cfar_cfarCore_cellUnderTest__T_15; // @[CFARUtils.scala 483:18]
  assign cfar_cfar_cfarCore_cellUnderTest_io_out_bits = cfar_cfar_cfarCore_cellUnderTest_cut; // @[CFARUtils.scala 481:18]
  assign cfar_cfar_cfarCore_cellUnderTest_io_lastOut = cfar_cfar_cfarCore_cellUnderTest_lastOut; // @[CFARUtils.scala 482:18]
  assign cfar_cfar_cfarCore_leadGuard__T_1 = cfar_cfar_cfarCore_leadGuard_io_in_ready & cfar_cfar_cfarCore_leadGuard_io_in_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_leadGuard__T_2 = cfar_cfar_cfarCore_leadGuard_last & cfar_cfar_cfarCore_leadGuard_io_out_ready; // @[CFARUtils.scala 385:34]
  assign cfar_cfar_cfarCore_leadGuard_en = cfar_cfar_cfarCore_leadGuard__T_1 | cfar_cfar_cfarCore_leadGuard__T_2; // @[CFARUtils.scala 385:25]
  assign cfar_cfar_cfarCore_leadGuard__T_3 = cfar_cfar_cfarCore_leadGuard_io_depth <= 4'h8; // @[CFARUtils.scala 345:18]
  assign cfar_cfar_cfarCore_leadGuard__T_5 = cfar_cfar_cfarCore_leadGuard__T_3 | cfar_cfar_cfarCore_leadGuard_reset; // @[CFARUtils.scala 345:11]
  assign cfar_cfar_cfarCore_leadGuard__T_6 = ~cfar_cfar_cfarCore_leadGuard__T_5; // @[CFARUtils.scala 345:11]
  assign cfar_cfar_cfarCore_leadGuard__T_8 = cfar_cfar_cfarCore_leadGuard_io_depth - 4'h1; // @[CFARUtils.scala 350:87]
  assign cfar_cfar_cfarCore_leadGuard__T_9 = 1'h1; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_13 = 4'h1 <= cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_14 = cfar_cfar_cfarCore_leadGuard__T_13; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_leadGuard__T_17 = 4'h2 <= cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_18 = cfar_cfar_cfarCore_leadGuard__T_17; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_leadGuard__T_21 = 4'h3 <= cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_22 = cfar_cfar_cfarCore_leadGuard__T_21; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_leadGuard__T_25 = 4'h4 <= cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_26 = cfar_cfar_cfarCore_leadGuard__T_25; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_leadGuard__T_29 = 4'h5 <= cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_30 = cfar_cfar_cfarCore_leadGuard__T_29; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_leadGuard__T_33 = 4'h6 <= cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_34 = cfar_cfar_cfarCore_leadGuard__T_33; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_leadGuard__T_37 = 4'h7 <= cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 350:78]
  assign cfar_cfar_cfarCore_leadGuard__T_38 = cfar_cfar_cfarCore_leadGuard__T_37; // @[CFARUtils.scala 350:94]
  assign cfar_cfar_cfarCore_leadGuard__T_39 = cfar_cfar_cfarCore_leadGuard__T_38 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_40 = cfar_cfar_cfarCore_leadGuard__T_34 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_41 = cfar_cfar_cfarCore_leadGuard__T_30 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_42 = cfar_cfar_cfarCore_leadGuard__T_26 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_43 = cfar_cfar_cfarCore_leadGuard__T_22 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_44 = cfar_cfar_cfarCore_leadGuard__T_18 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_45 = cfar_cfar_cfarCore_leadGuard__T_14 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_46 = cfar_cfar_cfarCore_leadGuard__T_9 & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_57 = cfar_cfar_cfarCore_leadGuard__T_8[2:0];
  assign cfar_cfar_cfarCore_leadGuard__T_59 = cfar_cfar_cfarCore_leadGuard_io_lastIn & cfar_cfar_cfarCore_leadGuard__T_1; // @[CFARUtils.scala 392:19]
  assign cfar_cfar_cfarCore_leadGuard__GEN_8 = cfar_cfar_cfarCore_leadGuard__T_59 | cfar_cfar_cfarCore_leadGuard_last; // @[CFARUtils.scala 392:36]
  assign cfar_cfar_cfarCore_leadGuard__T_62 = cfar_cfar_cfarCore_leadGuard_cntIn + 4'h1; // @[CFARUtils.scala 397:20]
  assign cfar_cfar_cfarCore_leadGuard__T_63 = cfar_cfar_cfarCore_leadGuard_io_depth > 4'h1; // @[CFARUtils.scala 400:18]
  assign cfar_cfar_cfarCore_leadGuard__T_66 = cfar_cfar_cfarCore_leadGuard_cntIn == cfar_cfar_cfarCore_leadGuard__T_8; // @[CFARUtils.scala 401:17]
  assign cfar_cfar_cfarCore_leadGuard__T_68 = cfar_cfar_cfarCore_leadGuard__T_66 & cfar_cfar_cfarCore_leadGuard__T_1; // @[CFARUtils.scala 401:36]
  assign cfar_cfar_cfarCore_leadGuard__GEN_10 = cfar_cfar_cfarCore_leadGuard__T_68 | cfar_cfar_cfarCore_leadGuard_InitialInDone; // @[CFARUtils.scala 401:53]
  assign cfar_cfar_cfarCore_leadGuard__T_70 = cfar_cfar_cfarCore_leadGuard_io_depth == 4'h1; // @[CFARUtils.scala 406:36]
  assign cfar_cfar_cfarCore_leadGuard__T_71 = cfar_cfar_cfarCore_leadGuard__T_1 & cfar_cfar_cfarCore_leadGuard__T_70; // @[CFARUtils.scala 406:24]
  assign cfar_cfar_cfarCore_leadGuard__GEN_11 = cfar_cfar_cfarCore_leadGuard__T_71 | cfar_cfar_cfarCore_leadGuard_InitialInDone; // @[CFARUtils.scala 406:45]
  assign cfar_cfar_cfarCore_leadGuard__T_73 = cfar_cfar_cfarCore_leadGuard_io_out_ready & cfar_cfar_cfarCore_leadGuard_io_out_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_leadGuard__T_112 = cfar_cfar_cfarCore_leadGuard__T_37 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_113 = cfar_cfar_cfarCore_leadGuard__T_33 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_114 = cfar_cfar_cfarCore_leadGuard__T_29 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_115 = cfar_cfar_cfarCore_leadGuard__T_25 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_116 = cfar_cfar_cfarCore_leadGuard__T_21 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_117 = cfar_cfar_cfarCore_leadGuard__T_17 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__T_118 = cfar_cfar_cfarCore_leadGuard__T_13 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadGuard__GEN_22 = 3'h1 == cfar_cfar_cfarCore_leadGuard__T_57 ? cfar_cfar_cfarCore_leadGuard__T_121 : cfar_cfar_cfarCore_leadGuard__T_120; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__GEN_23 = 3'h2 == cfar_cfar_cfarCore_leadGuard__T_57 ? cfar_cfar_cfarCore_leadGuard__T_122 : cfar_cfar_cfarCore_leadGuard__GEN_22; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__GEN_24 = 3'h3 == cfar_cfar_cfarCore_leadGuard__T_57 ? cfar_cfar_cfarCore_leadGuard__T_123 : cfar_cfar_cfarCore_leadGuard__GEN_23; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__GEN_25 = 3'h4 == cfar_cfar_cfarCore_leadGuard__T_57 ? cfar_cfar_cfarCore_leadGuard__T_124 : cfar_cfar_cfarCore_leadGuard__GEN_24; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__GEN_26 = 3'h5 == cfar_cfar_cfarCore_leadGuard__T_57 ? cfar_cfar_cfarCore_leadGuard__T_125 : cfar_cfar_cfarCore_leadGuard__GEN_25; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__GEN_27 = 3'h6 == cfar_cfar_cfarCore_leadGuard__T_57 ? cfar_cfar_cfarCore_leadGuard__T_126 : cfar_cfar_cfarCore_leadGuard__GEN_26; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__GEN_28 = 3'h7 == cfar_cfar_cfarCore_leadGuard__T_57 ? cfar_cfar_cfarCore_leadGuard__T_127 : cfar_cfar_cfarCore_leadGuard__GEN_27; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__T_132 = cfar_cfar_cfarCore_leadGuard__GEN_28 & cfar_cfar_cfarCore_leadGuard__T_73; // @[CFARUtils.scala 414:17]
  assign cfar_cfar_cfarCore_leadGuard__T_134 = ~cfar_cfar_cfarCore_leadGuard_InitialInDone; // @[CFARUtils.scala 420:36]
  assign cfar_cfar_cfarCore_leadGuard__T_136 = ~cfar_cfar_cfarCore_leadGuard_last; // @[CFARUtils.scala 421:36]
  assign cfar_cfar_cfarCore_leadGuard__T_138 = cfar_cfar_cfarCore_leadGuard_io_depth == 4'h0; // @[CFARUtils.scala 426:37]
  assign cfar_cfar_cfarCore_leadGuard__T_141 = cfar_cfar_cfarCore_leadGuard_io_out_ready & cfar_cfar_cfarCore_leadGuard__T_136; // @[CFARUtils.scala 426:91]
  assign cfar_cfar_cfarCore_leadGuard__T_142 = cfar_cfar_cfarCore_leadGuard__T_134 | cfar_cfar_cfarCore_leadGuard__T_141; // @[CFARUtils.scala 426:75]
  assign cfar_cfar_cfarCore_leadGuard__GEN_33 = 3'h1 == cfar_cfar_cfarCore_leadGuard__T_57 ? $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_1) : $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_0); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_leadGuard__GEN_34 = 3'h2 == cfar_cfar_cfarCore_leadGuard__T_57 ? $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_2) : $signed(cfar_cfar_cfarCore_leadGuard__GEN_33); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_leadGuard__GEN_35 = 3'h3 == cfar_cfar_cfarCore_leadGuard__T_57 ? $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_3) : $signed(cfar_cfar_cfarCore_leadGuard__GEN_34); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_leadGuard__GEN_36 = 3'h4 == cfar_cfar_cfarCore_leadGuard__T_57 ? $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_4) : $signed(cfar_cfar_cfarCore_leadGuard__GEN_35); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_leadGuard__GEN_37 = 3'h5 == cfar_cfar_cfarCore_leadGuard__T_57 ? $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_5) : $signed(cfar_cfar_cfarCore_leadGuard__GEN_36); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_leadGuard__GEN_38 = 3'h6 == cfar_cfar_cfarCore_leadGuard__T_57 ? $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_6) : $signed(cfar_cfar_cfarCore_leadGuard__GEN_37); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_leadGuard__GEN_39 = 3'h7 == cfar_cfar_cfarCore_leadGuard__T_57 ? $signed(cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_7) : $signed(cfar_cfar_cfarCore_leadGuard__GEN_38); // @[CFARUtils.scala 433:24]
  assign cfar_cfar_cfarCore_leadGuard__T_151 = cfar_cfar_cfarCore_leadGuard_InitialInDone & cfar_cfar_cfarCore_leadGuard_io_in_valid; // @[CFARUtils.scala 436:70]
  assign cfar_cfar_cfarCore_leadGuard__T_152 = cfar_cfar_cfarCore_leadGuard_last & cfar_cfar_cfarCore_leadGuard_en; // @[CFARUtils.scala 436:94]
  assign cfar_cfar_cfarCore_leadGuard__T_153 = cfar_cfar_cfarCore_leadGuard__T_151 | cfar_cfar_cfarCore_leadGuard__T_152; // @[CFARUtils.scala 436:85]
  assign cfar_cfar_cfarCore_leadGuard_io_in_ready = cfar_cfar_cfarCore_leadGuard__T_138 ? cfar_cfar_cfarCore_leadGuard_io_out_ready : cfar_cfar_cfarCore_leadGuard__T_142; // @[CFARUtils.scala 426:20]
  assign cfar_cfar_cfarCore_leadGuard_io_out_valid = cfar_cfar_cfarCore_leadGuard__T_138 ? cfar_cfar_cfarCore_leadGuard_io_in_valid : cfar_cfar_cfarCore_leadGuard__T_153; // @[CFARUtils.scala 436:18]
  assign cfar_cfar_cfarCore_leadGuard_io_out_bits = cfar_cfar_cfarCore_leadGuard__T_138 ? $signed(cfar_cfar_cfarCore_leadGuard_io_in_bits) : $signed(cfar_cfar_cfarCore_leadGuard__GEN_39); // @[CFARUtils.scala 433:18]
  assign cfar_cfar_cfarCore_leadGuard_io_lastOut = cfar_cfar_cfarCore_leadGuard__T_138 ? cfar_cfar_cfarCore_leadGuard__T_59 : cfar_cfar_cfarCore_leadGuard__GEN_28; // @[CFARUtils.scala 435:18]
  assign cfar_cfar_cfarCore_leadWindow_mem__T_423_addr = cfar_cfar_cfarCore_leadWindow_readIdx;
  assign cfar_cfar_cfarCore_leadWindow_mem__T_423_data = cfar_cfar_cfarCore_leadWindow_mem[cfar_cfar_cfarCore_leadWindow_mem__T_423_addr]; // @[CFARUtils.scala 505:26]
  assign cfar_cfar_cfarCore_leadWindow_mem__T_418_data = cfar_cfar_cfarCore_leadWindow_io_in_bits;
  assign cfar_cfar_cfarCore_leadWindow_mem__T_418_addr = cfar_cfar_cfarCore_leadWindow_writeIdxReg;
  assign cfar_cfar_cfarCore_leadWindow_mem__T_418_mask = 1'h1;
  assign cfar_cfar_cfarCore_leadWindow_mem__T_418_en = cfar_cfar_cfarCore_leadWindow_en & cfar_cfar_cfarCore_leadWindow__T_416;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_14_addr = 1'h0;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_14_data = cfar_cfar_cfarCore_leadWindow_outputQueue__T[cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_14_addr]; // @[Decoupled.scala 209:24]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_data = cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_bits;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_addr = 1'h0;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_mask = 1'h1;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_en = cfar_cfar_cfarCore_leadWindow_outputQueue__T_3 ? cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_7 : cfar_cfar_cfarCore_leadWindow_outputQueue__T_6;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T_3 = ~cfar_cfar_cfarCore_leadWindow_outputQueue__T_1; // @[Decoupled.scala 215:36]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T_6 = cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_ready & cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T_8 = cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_ready & cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_7 = cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_ready ? 1'h0 : cfar_cfar_cfarCore_leadWindow_outputQueue__T_6; // @[Decoupled.scala 240:27]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_10 = cfar_cfar_cfarCore_leadWindow_outputQueue__T_3 ? cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_7 : cfar_cfar_cfarCore_leadWindow_outputQueue__T_6; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_9 = cfar_cfar_cfarCore_leadWindow_outputQueue__T_3 ? 1'h0 : cfar_cfar_cfarCore_leadWindow_outputQueue__T_8; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T_11 = cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_10 != cfar_cfar_cfarCore_leadWindow_outputQueue__GEN_9; // @[Decoupled.scala 227:16]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue__T_12 = ~cfar_cfar_cfarCore_leadWindow_outputQueue__T_3; // @[Decoupled.scala 231:19]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_ready = cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_ready | cfar_cfar_cfarCore_leadWindow_outputQueue__T_3; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_valid = cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_valid | cfar_cfar_cfarCore_leadWindow_outputQueue__T_12; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_bits = cfar_cfar_cfarCore_leadWindow_outputQueue__T_3 ? $signed(cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_bits) : $signed(cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_14_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign cfar_cfar_cfarCore_leadWindow__T = cfar_cfar_cfarCore_leadWindow_io_in_ready & cfar_cfar_cfarCore_leadWindow_io_in_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_leadWindow__T_1 = cfar_cfar_cfarCore_leadWindow_last & cfar_cfar_cfarCore_leadWindow_io_out_ready; // @[CFARUtils.scala 511:45]
  assign cfar_cfar_cfarCore_leadWindow_en = cfar_cfar_cfarCore_leadWindow__T | cfar_cfar_cfarCore_leadWindow__T_1; // @[CFARUtils.scala 511:36]
  assign cfar_cfar_cfarCore_leadWindow__T_3 = cfar_cfar_cfarCore_leadWindow_writeIdxReg + 6'h1; // @[CFARUtils.scala 515:21]
  assign cfar_cfar_cfarCore_leadWindow__GEN_140 = {{1'd0}, cfar_cfar_cfarCore_leadWindow__T_3}; // @[CFARUtils.scala 515:27]
  assign cfar_cfar_cfarCore_leadWindow__T_4 = cfar_cfar_cfarCore_leadWindow__GEN_140 >= cfar_cfar_cfarCore_leadWindow_io_depth; // @[CFARUtils.scala 515:27]
  assign cfar_cfar_cfarCore_leadWindow__GEN_141 = {{1'd0}, cfar_cfar_cfarCore_leadWindow_writeIdxReg}; // @[CFARUtils.scala 516:28]
  assign cfar_cfar_cfarCore_leadWindow__T_6 = cfar_cfar_cfarCore_leadWindow__GEN_141 - cfar_cfar_cfarCore_leadWindow_io_depth; // @[CFARUtils.scala 516:28]
  assign cfar_cfar_cfarCore_leadWindow__T_8 = cfar_cfar_cfarCore_leadWindow__T_6 + 7'h1; // @[CFARUtils.scala 516:39]
  assign cfar_cfar_cfarCore_leadWindow__T_10 = 7'h40 + cfar_cfar_cfarCore_leadWindow__GEN_141; // @[CFARUtils.scala 518:27]
  assign cfar_cfar_cfarCore_leadWindow__T_12 = cfar_cfar_cfarCore_leadWindow__T_10 + 7'h1; // @[CFARUtils.scala 518:41]
  assign cfar_cfar_cfarCore_leadWindow__T_14 = cfar_cfar_cfarCore_leadWindow__T_12 - cfar_cfar_cfarCore_leadWindow_io_depth; // @[CFARUtils.scala 518:47]
  assign cfar_cfar_cfarCore_leadWindow__GEN_0 = cfar_cfar_cfarCore_leadWindow__T_4 ? cfar_cfar_cfarCore_leadWindow__T_8 : cfar_cfar_cfarCore_leadWindow__T_14; // @[CFARUtils.scala 515:40]
  assign cfar_cfar_cfarCore_leadWindow__T_16 = cfar_cfar_cfarCore_leadWindow_io_depth - 7'h1; // @[CFARUtils.scala 528:34]
  assign cfar_cfar_cfarCore_leadWindow__T_17 = cfar_cfar_cfarCore_leadWindow__GEN_141 == cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 528:21]
  assign cfar_cfar_cfarCore_leadWindow__T_19 = cfar_cfar_cfarCore_leadWindow__T_17 & cfar_cfar_cfarCore_leadWindow__T; // @[CFARUtils.scala 528:40]
  assign cfar_cfar_cfarCore_leadWindow__GEN_1 = cfar_cfar_cfarCore_leadWindow__T_19 | cfar_cfar_cfarCore_leadWindow_initialInDone; // @[CFARUtils.scala 528:57]
  assign cfar_cfar_cfarCore_leadWindow_fireLastIn = cfar_cfar_cfarCore_leadWindow_io_lastIn & cfar_cfar_cfarCore_leadWindow__T; // @[CFARUtils.scala 531:30]
  assign cfar_cfar_cfarCore_leadWindow__GEN_2 = cfar_cfar_cfarCore_leadWindow_fireLastIn | cfar_cfar_cfarCore_leadWindow_last; // @[CFARUtils.scala 533:21]
  assign cfar_cfar_cfarCore_leadWindow__T_21 = cfar_cfar_cfarCore_leadWindow_io_out_ready & cfar_cfar_cfarCore_leadWindow_io_out_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_leadWindow__T_22 = cfar_cfar_cfarCore_leadWindow_io_depth <= 7'h40; // @[CFARUtils.scala 330:18]
  assign cfar_cfar_cfarCore_leadWindow__T_24 = cfar_cfar_cfarCore_leadWindow__T_22 | cfar_cfar_cfarCore_leadWindow_reset; // @[CFARUtils.scala 330:11]
  assign cfar_cfar_cfarCore_leadWindow__T_25 = ~cfar_cfar_cfarCore_leadWindow__T_24; // @[CFARUtils.scala 330:11]
  assign cfar_cfar_cfarCore_leadWindow__T_33 = 7'h1 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_37 = 7'h2 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_41 = 7'h3 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_45 = 7'h4 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_49 = 7'h5 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_53 = 7'h6 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_57 = 7'h7 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_61 = 7'h8 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_65 = 7'h9 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_69 = 7'ha <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_73 = 7'hb <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_77 = 7'hc <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_81 = 7'hd <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_85 = 7'he <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_89 = 7'hf <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_93 = 7'h10 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_97 = 7'h11 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_101 = 7'h12 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_105 = 7'h13 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_109 = 7'h14 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_113 = 7'h15 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_117 = 7'h16 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_121 = 7'h17 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_125 = 7'h18 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_129 = 7'h19 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_133 = 7'h1a <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_137 = 7'h1b <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_141 = 7'h1c <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_145 = 7'h1d <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_149 = 7'h1e <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_153 = 7'h1f <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_157 = 7'h20 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_161 = 7'h21 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_165 = 7'h22 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_169 = 7'h23 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_173 = 7'h24 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_177 = 7'h25 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_181 = 7'h26 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_185 = 7'h27 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_189 = 7'h28 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_193 = 7'h29 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_197 = 7'h2a <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_201 = 7'h2b <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_205 = 7'h2c <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_209 = 7'h2d <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_213 = 7'h2e <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_217 = 7'h2f <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_221 = 7'h30 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_225 = 7'h31 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_229 = 7'h32 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_233 = 7'h33 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_237 = 7'h34 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_241 = 7'h35 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_245 = 7'h36 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_249 = 7'h37 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_253 = 7'h38 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_257 = 7'h39 <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_261 = 7'h3a <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_265 = 7'h3b <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_269 = 7'h3c <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_273 = 7'h3d <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_277 = 7'h3e <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_281 = 7'h3f <= cfar_cfar_cfarCore_leadWindow__T_16; // @[CFARUtils.scala 335:78]
  assign cfar_cfar_cfarCore_leadWindow__T_284 = cfar_cfar_cfarCore_leadWindow__T_281 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_285 = cfar_cfar_cfarCore_leadWindow__T_277 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_286 = cfar_cfar_cfarCore_leadWindow__T_273 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_287 = cfar_cfar_cfarCore_leadWindow__T_269 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_288 = cfar_cfar_cfarCore_leadWindow__T_265 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_289 = cfar_cfar_cfarCore_leadWindow__T_261 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_290 = cfar_cfar_cfarCore_leadWindow__T_257 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_291 = cfar_cfar_cfarCore_leadWindow__T_253 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_292 = cfar_cfar_cfarCore_leadWindow__T_249 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_293 = cfar_cfar_cfarCore_leadWindow__T_245 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_294 = cfar_cfar_cfarCore_leadWindow__T_241 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_295 = cfar_cfar_cfarCore_leadWindow__T_237 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_296 = cfar_cfar_cfarCore_leadWindow__T_233 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_297 = cfar_cfar_cfarCore_leadWindow__T_229 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_298 = cfar_cfar_cfarCore_leadWindow__T_225 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_299 = cfar_cfar_cfarCore_leadWindow__T_221 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_300 = cfar_cfar_cfarCore_leadWindow__T_217 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_301 = cfar_cfar_cfarCore_leadWindow__T_213 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_302 = cfar_cfar_cfarCore_leadWindow__T_209 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_303 = cfar_cfar_cfarCore_leadWindow__T_205 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_304 = cfar_cfar_cfarCore_leadWindow__T_201 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_305 = cfar_cfar_cfarCore_leadWindow__T_197 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_306 = cfar_cfar_cfarCore_leadWindow__T_193 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_307 = cfar_cfar_cfarCore_leadWindow__T_189 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_308 = cfar_cfar_cfarCore_leadWindow__T_185 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_309 = cfar_cfar_cfarCore_leadWindow__T_181 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_310 = cfar_cfar_cfarCore_leadWindow__T_177 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_311 = cfar_cfar_cfarCore_leadWindow__T_173 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_312 = cfar_cfar_cfarCore_leadWindow__T_169 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_313 = cfar_cfar_cfarCore_leadWindow__T_165 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_314 = cfar_cfar_cfarCore_leadWindow__T_161 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_315 = cfar_cfar_cfarCore_leadWindow__T_157 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_316 = cfar_cfar_cfarCore_leadWindow__T_153 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_317 = cfar_cfar_cfarCore_leadWindow__T_149 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_318 = cfar_cfar_cfarCore_leadWindow__T_145 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_319 = cfar_cfar_cfarCore_leadWindow__T_141 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_320 = cfar_cfar_cfarCore_leadWindow__T_137 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_321 = cfar_cfar_cfarCore_leadWindow__T_133 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_322 = cfar_cfar_cfarCore_leadWindow__T_129 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_323 = cfar_cfar_cfarCore_leadWindow__T_125 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_324 = cfar_cfar_cfarCore_leadWindow__T_121 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_325 = cfar_cfar_cfarCore_leadWindow__T_117 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_326 = cfar_cfar_cfarCore_leadWindow__T_113 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_327 = cfar_cfar_cfarCore_leadWindow__T_109 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_328 = cfar_cfar_cfarCore_leadWindow__T_105 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_329 = cfar_cfar_cfarCore_leadWindow__T_101 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_330 = cfar_cfar_cfarCore_leadWindow__T_97 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_331 = cfar_cfar_cfarCore_leadWindow__T_93 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_332 = cfar_cfar_cfarCore_leadWindow__T_89 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_333 = cfar_cfar_cfarCore_leadWindow__T_85 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_334 = cfar_cfar_cfarCore_leadWindow__T_81 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_335 = cfar_cfar_cfarCore_leadWindow__T_77 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_336 = cfar_cfar_cfarCore_leadWindow__T_73 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_337 = cfar_cfar_cfarCore_leadWindow__T_69 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_338 = cfar_cfar_cfarCore_leadWindow__T_65 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_339 = cfar_cfar_cfarCore_leadWindow__T_61 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_340 = cfar_cfar_cfarCore_leadWindow__T_57 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_341 = cfar_cfar_cfarCore_leadWindow__T_53 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_342 = cfar_cfar_cfarCore_leadWindow__T_49 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_343 = cfar_cfar_cfarCore_leadWindow__T_45 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_344 = cfar_cfar_cfarCore_leadWindow__T_41 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_345 = cfar_cfar_cfarCore_leadWindow__T_37 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_346 = cfar_cfar_cfarCore_leadWindow__T_33 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 319:37]
  assign cfar_cfar_cfarCore_leadWindow__T_414 = cfar_cfar_cfarCore_leadWindow__T_16[5:0];
  assign cfar_cfar_cfarCore_leadWindow__GEN_68 = 6'h1 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_349 : cfar_cfar_cfarCore_leadWindow__T_348; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_69 = 6'h2 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_350 : cfar_cfar_cfarCore_leadWindow__GEN_68; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_70 = 6'h3 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_351 : cfar_cfar_cfarCore_leadWindow__GEN_69; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_71 = 6'h4 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_352 : cfar_cfar_cfarCore_leadWindow__GEN_70; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_72 = 6'h5 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_353 : cfar_cfar_cfarCore_leadWindow__GEN_71; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_73 = 6'h6 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_354 : cfar_cfar_cfarCore_leadWindow__GEN_72; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_74 = 6'h7 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_355 : cfar_cfar_cfarCore_leadWindow__GEN_73; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_75 = 6'h8 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_356 : cfar_cfar_cfarCore_leadWindow__GEN_74; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_76 = 6'h9 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_357 : cfar_cfar_cfarCore_leadWindow__GEN_75; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_77 = 6'ha == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_358 : cfar_cfar_cfarCore_leadWindow__GEN_76; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_78 = 6'hb == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_359 : cfar_cfar_cfarCore_leadWindow__GEN_77; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_79 = 6'hc == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_360 : cfar_cfar_cfarCore_leadWindow__GEN_78; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_80 = 6'hd == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_361 : cfar_cfar_cfarCore_leadWindow__GEN_79; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_81 = 6'he == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_362 : cfar_cfar_cfarCore_leadWindow__GEN_80; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_82 = 6'hf == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_363 : cfar_cfar_cfarCore_leadWindow__GEN_81; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_83 = 6'h10 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_364 : cfar_cfar_cfarCore_leadWindow__GEN_82; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_84 = 6'h11 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_365 : cfar_cfar_cfarCore_leadWindow__GEN_83; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_85 = 6'h12 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_366 : cfar_cfar_cfarCore_leadWindow__GEN_84; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_86 = 6'h13 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_367 : cfar_cfar_cfarCore_leadWindow__GEN_85; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_87 = 6'h14 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_368 : cfar_cfar_cfarCore_leadWindow__GEN_86; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_88 = 6'h15 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_369 : cfar_cfar_cfarCore_leadWindow__GEN_87; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_89 = 6'h16 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_370 : cfar_cfar_cfarCore_leadWindow__GEN_88; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_90 = 6'h17 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_371 : cfar_cfar_cfarCore_leadWindow__GEN_89; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_91 = 6'h18 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_372 : cfar_cfar_cfarCore_leadWindow__GEN_90; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_92 = 6'h19 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_373 : cfar_cfar_cfarCore_leadWindow__GEN_91; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_93 = 6'h1a == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_374 : cfar_cfar_cfarCore_leadWindow__GEN_92; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_94 = 6'h1b == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_375 : cfar_cfar_cfarCore_leadWindow__GEN_93; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_95 = 6'h1c == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_376 : cfar_cfar_cfarCore_leadWindow__GEN_94; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_96 = 6'h1d == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_377 : cfar_cfar_cfarCore_leadWindow__GEN_95; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_97 = 6'h1e == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_378 : cfar_cfar_cfarCore_leadWindow__GEN_96; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_98 = 6'h1f == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_379 : cfar_cfar_cfarCore_leadWindow__GEN_97; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_99 = 6'h20 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_380 : cfar_cfar_cfarCore_leadWindow__GEN_98; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_100 = 6'h21 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_381 : cfar_cfar_cfarCore_leadWindow__GEN_99; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_101 = 6'h22 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_382 : cfar_cfar_cfarCore_leadWindow__GEN_100; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_102 = 6'h23 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_383 : cfar_cfar_cfarCore_leadWindow__GEN_101; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_103 = 6'h24 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_384 : cfar_cfar_cfarCore_leadWindow__GEN_102; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_104 = 6'h25 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_385 : cfar_cfar_cfarCore_leadWindow__GEN_103; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_105 = 6'h26 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_386 : cfar_cfar_cfarCore_leadWindow__GEN_104; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_106 = 6'h27 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_387 : cfar_cfar_cfarCore_leadWindow__GEN_105; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_107 = 6'h28 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_388 : cfar_cfar_cfarCore_leadWindow__GEN_106; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_108 = 6'h29 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_389 : cfar_cfar_cfarCore_leadWindow__GEN_107; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_109 = 6'h2a == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_390 : cfar_cfar_cfarCore_leadWindow__GEN_108; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_110 = 6'h2b == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_391 : cfar_cfar_cfarCore_leadWindow__GEN_109; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_111 = 6'h2c == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_392 : cfar_cfar_cfarCore_leadWindow__GEN_110; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_112 = 6'h2d == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_393 : cfar_cfar_cfarCore_leadWindow__GEN_111; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_113 = 6'h2e == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_394 : cfar_cfar_cfarCore_leadWindow__GEN_112; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_114 = 6'h2f == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_395 : cfar_cfar_cfarCore_leadWindow__GEN_113; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_115 = 6'h30 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_396 : cfar_cfar_cfarCore_leadWindow__GEN_114; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_116 = 6'h31 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_397 : cfar_cfar_cfarCore_leadWindow__GEN_115; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_117 = 6'h32 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_398 : cfar_cfar_cfarCore_leadWindow__GEN_116; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_118 = 6'h33 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_399 : cfar_cfar_cfarCore_leadWindow__GEN_117; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_119 = 6'h34 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_400 : cfar_cfar_cfarCore_leadWindow__GEN_118; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_120 = 6'h35 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_401 : cfar_cfar_cfarCore_leadWindow__GEN_119; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_121 = 6'h36 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_402 : cfar_cfar_cfarCore_leadWindow__GEN_120; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_122 = 6'h37 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_403 : cfar_cfar_cfarCore_leadWindow__GEN_121; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_123 = 6'h38 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_404 : cfar_cfar_cfarCore_leadWindow__GEN_122; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_124 = 6'h39 == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_405 : cfar_cfar_cfarCore_leadWindow__GEN_123; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_125 = 6'h3a == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_406 : cfar_cfar_cfarCore_leadWindow__GEN_124; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_126 = 6'h3b == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_407 : cfar_cfar_cfarCore_leadWindow__GEN_125; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_127 = 6'h3c == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_408 : cfar_cfar_cfarCore_leadWindow__GEN_126; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_128 = 6'h3d == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_409 : cfar_cfar_cfarCore_leadWindow__GEN_127; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_129 = 6'h3e == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_410 : cfar_cfar_cfarCore_leadWindow__GEN_128; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__GEN_130 = 6'h3f == cfar_cfar_cfarCore_leadWindow__T_414 ? cfar_cfar_cfarCore_leadWindow__T_411 : cfar_cfar_cfarCore_leadWindow__GEN_129; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow_resetAll = cfar_cfar_cfarCore_leadWindow__GEN_130 & cfar_cfar_cfarCore_leadWindow__T_21; // @[CFARUtils.scala 537:26]
  assign cfar_cfar_cfarCore_leadWindow__T_416 = ~cfar_cfar_cfarCore_leadWindow_resetAll; // @[CFARUtils.scala 544:15]
  assign cfar_cfar_cfarCore_leadWindow__T_417 = cfar_cfar_cfarCore_leadWindow_en & cfar_cfar_cfarCore_leadWindow__T_416; // @[CFARUtils.scala 544:12]
  assign cfar_cfar_cfarCore_leadWindow__T_419 = cfar_cfar_cfarCore_leadWindow_writeIdxReg < 6'h3f; // @[CFARUtils.scala 546:36]
  assign cfar_cfar_cfarCore_leadWindow__T_430 = cfar_cfar_cfarCore_leadWindow_writeIdxReg == 6'h0; // @[CFARUtils.scala 554:31]
  assign cfar_cfar_cfarCore_leadWindow__T_431 = ~cfar_cfar_cfarCore_leadWindow_initialInDone; // @[CFARUtils.scala 554:42]
  assign cfar_cfar_cfarCore_leadWindow__T_433 = ~cfar_cfar_cfarCore_leadWindow_last; // @[CFARUtils.scala 555:36]
  assign cfar_cfar_cfarCore_leadWindow__T_437 = cfar_cfar_cfarCore_leadWindow_initialInDone & cfar_cfar_cfarCore_leadWindow_io_in_valid; // @[CFARUtils.scala 568:33]
  assign cfar_cfar_cfarCore_leadWindow__T_438 = cfar_cfar_cfarCore_leadWindow_last & cfar_cfar_cfarCore_leadWindow_en; // @[CFARUtils.scala 568:57]
  assign cfar_cfar_cfarCore_leadWindow_readIdx = cfar_cfar_cfarCore_leadWindow__GEN_0[5:0]; // @[CFARUtils.scala 506:27 CFARUtils.scala 516:13 CFARUtils.scala 518:13]
  assign cfar_cfar_cfarCore_leadWindow_io_in_ready = cfar_cfar_cfarCore_leadWindow_io_out_ready & cfar_cfar_cfarCore_leadWindow__T_433; // @[CFARUtils.scala 562:18]
  assign cfar_cfar_cfarCore_leadWindow_io_out_valid = cfar_cfar_cfarCore_leadWindow__T_437 | cfar_cfar_cfarCore_leadWindow__T_438; // @[CFARUtils.scala 568:16]
  assign cfar_cfar_cfarCore_leadWindow_io_out_bits = cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_bits; // @[CFARUtils.scala 565:16]
  assign cfar_cfar_cfarCore_leadWindow_io_memFull = cfar_cfar_cfarCore_leadWindow_initialInDone & cfar_cfar_cfarCore_leadWindow__T_433; // @[CFARUtils.scala 555:16]
  assign cfar_cfar_cfarCore_leadWindow_io_memEmpty = cfar_cfar_cfarCore_leadWindow__T_430 & cfar_cfar_cfarCore_leadWindow__T_431; // @[CFARUtils.scala 554:16]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_clock = cfar_cfar_cfarCore_leadWindow_clock;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_reset = cfar_cfar_cfarCore_leadWindow_reset;
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_valid = cfar_cfar_cfarCore_leadWindow_validPrev; // @[CFARUtils.scala 550:28]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_io_enq_bits = cfar_cfar_cfarCore_leadWindow__T_426; // @[CFARUtils.scala 551:27]
  assign cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_ready = cfar_cfar_cfarCore_leadWindow__T | cfar_cfar_cfarCore_leadWindow__T_1; // @[CFARUtils.scala 552:28]
  assign cfar_cfar_cfarCore_Queue__T_peak__T_18_addr = cfar_cfar_cfarCore_Queue_value_1;
  assign cfar_cfar_cfarCore_Queue__T_peak__T_18_data = cfar_cfar_cfarCore_Queue__T_peak[cfar_cfar_cfarCore_Queue__T_peak__T_18_addr]; // @[Decoupled.scala 209:24]
  assign cfar_cfar_cfarCore_Queue__T_peak__T_10_data = cfar_cfar_cfarCore_Queue_io_enq_bits_peak;
  assign cfar_cfar_cfarCore_Queue__T_peak__T_10_addr = cfar_cfar_cfarCore_Queue_value;
  assign cfar_cfar_cfarCore_Queue__T_peak__T_10_mask = 1'h1;
  assign cfar_cfar_cfarCore_Queue__T_peak__T_10_en = cfar_cfar_cfarCore_Queue__T_4 ? cfar_cfar_cfarCore_Queue__GEN_11 : cfar_cfar_cfarCore_Queue__T_6;
  assign cfar_cfar_cfarCore_Queue__T_cut__T_18_addr = cfar_cfar_cfarCore_Queue_value_1;
  assign cfar_cfar_cfarCore_Queue__T_cut__T_18_data = cfar_cfar_cfarCore_Queue__T_cut[cfar_cfar_cfarCore_Queue__T_cut__T_18_addr]; // @[Decoupled.scala 209:24]
  assign cfar_cfar_cfarCore_Queue__T_cut__T_10_data = cfar_cfar_cfarCore_Queue_io_enq_bits_cut;
  assign cfar_cfar_cfarCore_Queue__T_cut__T_10_addr = cfar_cfar_cfarCore_Queue_value;
  assign cfar_cfar_cfarCore_Queue__T_cut__T_10_mask = 1'h1;
  assign cfar_cfar_cfarCore_Queue__T_cut__T_10_en = cfar_cfar_cfarCore_Queue__T_4 ? cfar_cfar_cfarCore_Queue__GEN_11 : cfar_cfar_cfarCore_Queue__T_6;
  assign cfar_cfar_cfarCore_Queue__T_threshold__T_18_addr = cfar_cfar_cfarCore_Queue_value_1;
  assign cfar_cfar_cfarCore_Queue__T_threshold__T_18_data = cfar_cfar_cfarCore_Queue__T_threshold[cfar_cfar_cfarCore_Queue__T_threshold__T_18_addr]; // @[Decoupled.scala 209:24]
  assign cfar_cfar_cfarCore_Queue__T_threshold__T_10_data = cfar_cfar_cfarCore_Queue_io_enq_bits_threshold;
  assign cfar_cfar_cfarCore_Queue__T_threshold__T_10_addr = cfar_cfar_cfarCore_Queue_value;
  assign cfar_cfar_cfarCore_Queue__T_threshold__T_10_mask = 1'h1;
  assign cfar_cfar_cfarCore_Queue__T_threshold__T_10_en = cfar_cfar_cfarCore_Queue__T_4 ? cfar_cfar_cfarCore_Queue__GEN_11 : cfar_cfar_cfarCore_Queue__T_6;
  assign cfar_cfar_cfarCore_Queue__T_2 = cfar_cfar_cfarCore_Queue_value == cfar_cfar_cfarCore_Queue_value_1; // @[Decoupled.scala 214:41]
  assign cfar_cfar_cfarCore_Queue__T_3 = ~cfar_cfar_cfarCore_Queue__T_1; // @[Decoupled.scala 215:36]
  assign cfar_cfar_cfarCore_Queue__T_4 = cfar_cfar_cfarCore_Queue__T_2 & cfar_cfar_cfarCore_Queue__T_3; // @[Decoupled.scala 215:33]
  assign cfar_cfar_cfarCore_Queue__T_5 = cfar_cfar_cfarCore_Queue__T_2 & cfar_cfar_cfarCore_Queue__T_1; // @[Decoupled.scala 216:32]
  assign cfar_cfar_cfarCore_Queue__T_6 = cfar_cfar_cfarCore_Queue_io_enq_ready & cfar_cfar_cfarCore_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_Queue__T_8 = cfar_cfar_cfarCore_Queue_io_deq_ready & cfar_cfar_cfarCore_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_Queue__T_12 = cfar_cfar_cfarCore_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign cfar_cfar_cfarCore_Queue__GEN_11 = cfar_cfar_cfarCore_Queue_io_deq_ready ? 1'h0 : cfar_cfar_cfarCore_Queue__T_6; // @[Decoupled.scala 240:27]
  assign cfar_cfar_cfarCore_Queue__GEN_16 = cfar_cfar_cfarCore_Queue__T_4 ? cfar_cfar_cfarCore_Queue__GEN_11 : cfar_cfar_cfarCore_Queue__T_6; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_Queue__T_14 = cfar_cfar_cfarCore_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign cfar_cfar_cfarCore_Queue__GEN_15 = cfar_cfar_cfarCore_Queue__T_4 ? 1'h0 : cfar_cfar_cfarCore_Queue__T_8; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_Queue__T_15 = cfar_cfar_cfarCore_Queue__GEN_16 != cfar_cfar_cfarCore_Queue__GEN_15; // @[Decoupled.scala 227:16]
  assign cfar_cfar_cfarCore_Queue__T_16 = ~cfar_cfar_cfarCore_Queue__T_4; // @[Decoupled.scala 231:19]
  assign cfar_cfar_cfarCore_Queue_io_enq_ready = ~cfar_cfar_cfarCore_Queue__T_5; // @[Decoupled.scala 232:16]
  assign cfar_cfar_cfarCore_Queue_io_deq_valid = cfar_cfar_cfarCore_Queue_io_enq_valid | cfar_cfar_cfarCore_Queue__T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign cfar_cfar_cfarCore_Queue_io_deq_bits_peak = cfar_cfar_cfarCore_Queue__T_4 ? cfar_cfar_cfarCore_Queue_io_enq_bits_peak : cfar_cfar_cfarCore_Queue__T_peak__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign cfar_cfar_cfarCore_Queue_io_deq_bits_cut = cfar_cfar_cfarCore_Queue__T_4 ? $signed(cfar_cfar_cfarCore_Queue_io_enq_bits_cut) : $signed(cfar_cfar_cfarCore_Queue__T_cut__T_18_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign cfar_cfar_cfarCore_Queue_io_deq_bits_threshold = cfar_cfar_cfarCore_Queue__T_4 ? $signed(cfar_cfar_cfarCore_Queue_io_enq_bits_threshold) : $signed(cfar_cfar_cfarCore_Queue__T_threshold__T_18_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign cfar_cfar_cfarCore_Queue_2__T__T_18_addr = cfar_cfar_cfarCore_Queue_2_value_1;
  assign cfar_cfar_cfarCore_Queue_2__T__T_18_data = cfar_cfar_cfarCore_Queue_2__T[cfar_cfar_cfarCore_Queue_2__T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign cfar_cfar_cfarCore_Queue_2__T__T_10_data = cfar_cfar_cfarCore_Queue_2_io_enq_bits;
  assign cfar_cfar_cfarCore_Queue_2__T__T_10_addr = cfar_cfar_cfarCore_Queue_2_value;
  assign cfar_cfar_cfarCore_Queue_2__T__T_10_mask = 1'h1;
  assign cfar_cfar_cfarCore_Queue_2__T__T_10_en = cfar_cfar_cfarCore_Queue_2__T_4 ? cfar_cfar_cfarCore_Queue_2__GEN_9 : cfar_cfar_cfarCore_Queue_2__T_6;
  assign cfar_cfar_cfarCore_Queue_2__T_2 = cfar_cfar_cfarCore_Queue_2_value == cfar_cfar_cfarCore_Queue_2_value_1; // @[Decoupled.scala 214:41]
  assign cfar_cfar_cfarCore_Queue_2__T_3 = ~cfar_cfar_cfarCore_Queue_2__T_1; // @[Decoupled.scala 215:36]
  assign cfar_cfar_cfarCore_Queue_2__T_4 = cfar_cfar_cfarCore_Queue_2__T_2 & cfar_cfar_cfarCore_Queue_2__T_3; // @[Decoupled.scala 215:33]
  assign cfar_cfar_cfarCore_Queue_2__T_5 = cfar_cfar_cfarCore_Queue_2__T_2 & cfar_cfar_cfarCore_Queue_2__T_1; // @[Decoupled.scala 216:32]
  assign cfar_cfar_cfarCore_Queue_2__T_6 = cfar_cfar_cfarCore_Queue_2_io_enq_ready & cfar_cfar_cfarCore_Queue_2_io_enq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_Queue_2__T_8 = cfar_cfar_cfarCore_Queue_2_io_deq_ready & cfar_cfar_cfarCore_Queue_2_io_deq_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore_Queue_2__T_12 = cfar_cfar_cfarCore_Queue_2_value + 1'h1; // @[Counter.scala 39:22]
  assign cfar_cfar_cfarCore_Queue_2__GEN_9 = cfar_cfar_cfarCore_Queue_2_io_deq_ready ? 1'h0 : cfar_cfar_cfarCore_Queue_2__T_6; // @[Decoupled.scala 240:27]
  assign cfar_cfar_cfarCore_Queue_2__GEN_12 = cfar_cfar_cfarCore_Queue_2__T_4 ? cfar_cfar_cfarCore_Queue_2__GEN_9 : cfar_cfar_cfarCore_Queue_2__T_6; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_Queue_2__T_14 = cfar_cfar_cfarCore_Queue_2_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign cfar_cfar_cfarCore_Queue_2__GEN_11 = cfar_cfar_cfarCore_Queue_2__T_4 ? 1'h0 : cfar_cfar_cfarCore_Queue_2__T_8; // @[Decoupled.scala 237:18]
  assign cfar_cfar_cfarCore_Queue_2__T_15 = cfar_cfar_cfarCore_Queue_2__GEN_12 != cfar_cfar_cfarCore_Queue_2__GEN_11; // @[Decoupled.scala 227:16]
  assign cfar_cfar_cfarCore_Queue_2__T_16 = ~cfar_cfar_cfarCore_Queue_2__T_4; // @[Decoupled.scala 231:19]
  assign cfar_cfar_cfarCore_Queue_2_io_enq_ready = ~cfar_cfar_cfarCore_Queue_2__T_5; // @[Decoupled.scala 232:16]
  assign cfar_cfar_cfarCore_Queue_2_io_deq_valid = cfar_cfar_cfarCore_Queue_2_io_enq_valid | cfar_cfar_cfarCore_Queue_2__T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign cfar_cfar_cfarCore_Queue_2_io_deq_bits = cfar_cfar_cfarCore_Queue_2__T_4 ? cfar_cfar_cfarCore_Queue_2_io_enq_bits : cfar_cfar_cfarCore_Queue_2__T__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign cfar_cfar_cfarCore__GEN_41 = {{3'd0}, cfar_cfar_cfarCore_io_guardCells}; // @[CFARCoreWithMem.scala 32:32]
  assign cfar_cfar_cfarCore__T = cfar_cfar_cfarCore_io_windowCells + cfar_cfar_cfarCore__GEN_41; // @[CFARCoreWithMem.scala 32:32]
  assign cfar_cfar_cfarCore_latency = cfar_cfar_cfarCore__T + 8'h1; // @[CFARCoreWithMem.scala 32:49]
  assign cfar_cfar_cfarCore__T_1 = 7'h2 * cfar_cfar_cfarCore_io_windowCells; // @[CFARCoreWithMem.scala 33:26]
  assign cfar_cfar_cfarCore__T_2 = 4'h2 * cfar_cfar_cfarCore_io_guardCells; // @[CFARCoreWithMem.scala 33:49]
  assign cfar_cfar_cfarCore__GEN_42 = {{3'd0}, cfar_cfar_cfarCore__T_2}; // @[CFARCoreWithMem.scala 33:43]
  assign cfar_cfar_cfarCore__T_4 = cfar_cfar_cfarCore__T_1 + cfar_cfar_cfarCore__GEN_42; // @[CFARCoreWithMem.scala 33:43]
  assign cfar_cfar_cfarCore__T_6 = cfar_cfar_cfarCore__T_4 + 9'h1; // @[CFARCoreWithMem.scala 33:65]
  assign cfar_cfar_cfarCore__GEN_43 = {{1'd0}, cfar_cfar_cfarCore__T_6}; // @[CFARCoreWithMem.scala 33:20]
  assign cfar_cfar_cfarCore__T_7 = cfar_cfar_cfarCore_io_fftWin > cfar_cfar_cfarCore__GEN_43; // @[CFARCoreWithMem.scala 33:20]
  assign cfar_cfar_cfarCore__T_9 = cfar_cfar_cfarCore__T_7 | cfar_cfar_cfarCore_reset; // @[CFARCoreWithMem.scala 33:9]
  assign cfar_cfar_cfarCore__T_10 = ~cfar_cfar_cfarCore__T_9; // @[CFARCoreWithMem.scala 33:9]
  assign cfar_cfar_cfarCore__T_11 = cfar_cfar_cfarCore_io_guardCells > 4'h0; // @[CFARCoreWithMem.scala 34:24]
  assign cfar_cfar_cfarCore__T_13 = cfar_cfar_cfarCore__T_11 | cfar_cfar_cfarCore_reset; // @[CFARCoreWithMem.scala 34:9]
  assign cfar_cfar_cfarCore__T_14 = ~cfar_cfar_cfarCore__T_13; // @[CFARCoreWithMem.scala 34:9]
  assign cfar_cfar_cfarCore__T_21 = cfar_cfar_cfarCore_io_in_ready & cfar_cfar_cfarCore_io_in_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore__T_23 = cfar_cfar_cfarCore_cntIn + 9'h1; // @[CFARCoreWithMem.scala 75:20]
  assign cfar_cfar_cfarCore__T_25 = cfar_cfar_cfarCore_latency - 9'h1; // @[CFARCoreWithMem.scala 77:28]
  assign cfar_cfar_cfarCore__T_26 = cfar_cfar_cfarCore_cntIn == cfar_cfar_cfarCore__T_25; // @[CFARCoreWithMem.scala 77:15]
  assign cfar_cfar_cfarCore__T_28 = cfar_cfar_cfarCore__T_26 & cfar_cfar_cfarCore__T_21; // @[CFARCoreWithMem.scala 77:35]
  assign cfar_cfar_cfarCore__GEN_2 = cfar_cfar_cfarCore__T_28 | cfar_cfar_cfarCore_initialInDone; // @[CFARCoreWithMem.scala 77:52]
  assign cfar_cfar_cfarCore__T_29 = cfar_cfar_cfarCore_io_out_ready & cfar_cfar_cfarCore_io_out_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore__T_30 = cfar_cfar_cfarCore_io_lastOut & cfar_cfar_cfarCore__T_29; // @[CFARCoreWithMem.scala 81:20]
  assign cfar_cfar_cfarCore__T_33 = cfar_cfar_cfarCore_cntOut + 9'h1; // @[CFARCoreWithMem.scala 85:22]
  assign cfar_cfar_cfarCore__T_35 = cfar_cfar_cfarCore_io_fftWin - 10'h1; // @[CFARCoreWithMem.scala 87:31]
  assign cfar_cfar_cfarCore__GEN_44 = {{1'd0}, cfar_cfar_cfarCore_cntOut}; // @[CFARCoreWithMem.scala 87:16]
  assign cfar_cfar_cfarCore__T_36 = cfar_cfar_cfarCore__GEN_44 == cfar_cfar_cfarCore__T_35; // @[CFARCoreWithMem.scala 87:16]
  assign cfar_cfar_cfarCore__T_38 = cfar_cfar_cfarCore__T_36 & cfar_cfar_cfarCore__T_29; // @[CFARCoreWithMem.scala 87:38]
  assign cfar_cfar_cfarCore__T_41 = cfar_cfar_cfarCore__T_38 | cfar_cfar_cfarCore__T_30; // @[CFARCoreWithMem.scala 87:55]
  assign cfar_cfar_cfarCore__T_42 = cfar_cfar_cfarCore_io_lastIn & cfar_cfar_cfarCore_io_in_valid; // @[CFARCoreWithMem.scala 93:19]
  assign cfar_cfar_cfarCore__GEN_6 = cfar_cfar_cfarCore__T_42 | cfar_cfar_cfarCore_flushing; // @[CFARCoreWithMem.scala 93:35]
  assign cfar_cfar_cfarCore__GEN_9 = cfar_cfar_cfarCore_io_lastOut | cfar_cfar_cfarCore_lastCut; // @[CFARCoreWithMem.scala 101:21]
  assign cfar_cfar_cfarCore__T_43 = cfar_cfar_cfarCore_leadWindow_io_memEmpty; // @[CFARCoreWithMem.scala 106:32]
  assign cfar_cfar_cfarCore__T_47 = cfar_cfar_cfarCore_laggWindow_io_out_ready & cfar_cfar_cfarCore_laggWindow_io_out_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore__GEN_45 = {{4{cfar_cfar_cfarCore_laggWindow_io_in_bits[15]}},cfar_cfar_cfarCore_laggWindow_io_in_bits}; // @[FixedPointTypeClass.scala 20:58]
  assign cfar_cfar_cfarCore__T_50 = $signed(cfar_cfar_cfarCore_sumlagg) + $signed(cfar_cfar_cfarCore__GEN_45); // @[FixedPointTypeClass.scala 20:58]
  assign cfar_cfar_cfarCore__GEN_46 = {{4{cfar_cfar_cfarCore_laggWindow_io_out_bits[15]}},cfar_cfar_cfarCore_laggWindow_io_out_bits}; // @[FixedPointTypeClass.scala 30:68]
  assign cfar_cfar_cfarCore__T_53 = $signed(cfar_cfar_cfarCore__T_50) - $signed(cfar_cfar_cfarCore__GEN_46); // @[FixedPointTypeClass.scala 30:68]
  assign cfar_cfar_cfarCore__T_59 = cfar_cfar_cfarCore_leadWindow_io_in_ready & cfar_cfar_cfarCore_leadWindow_io_in_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore__T_60 = cfar_cfar_cfarCore_leadWindow_io_out_ready & cfar_cfar_cfarCore_leadWindow_io_out_valid; // @[Decoupled.scala 40:37]
  assign cfar_cfar_cfarCore__GEN_48 = {{4{cfar_cfar_cfarCore_leadWindow_io_in_bits[15]}},cfar_cfar_cfarCore_leadWindow_io_in_bits}; // @[FixedPointTypeClass.scala 20:58]
  assign cfar_cfar_cfarCore__T_63 = $signed(cfar_cfar_cfarCore_sumlead) + $signed(cfar_cfar_cfarCore__GEN_48); // @[FixedPointTypeClass.scala 20:58]
  assign cfar_cfar_cfarCore__GEN_49 = {{4{cfar_cfar_cfarCore_leadWindow_io_out_bits[15]}},cfar_cfar_cfarCore_leadWindow_io_out_bits}; // @[FixedPointTypeClass.scala 30:68]
  assign cfar_cfar_cfarCore__T_66 = $signed(cfar_cfar_cfarCore__T_63) - $signed(cfar_cfar_cfarCore__GEN_49); // @[FixedPointTypeClass.scala 30:68]
  assign cfar_cfar_cfarCore_leftThr = $signed(cfar_cfar_cfarCore_sumlagg) >>> cfar_cfar_cfarCore_io_divSum; // @[FixedPointTypeClass.scala 118:51]
  assign cfar_cfar_cfarCore_rightThr = $signed(cfar_cfar_cfarCore_sumlead) >>> cfar_cfar_cfarCore_io_divSum; // @[FixedPointTypeClass.scala 118:51]
  assign cfar_cfar_cfarCore__T_70 = $signed(cfar_cfar_cfarCore_leftThr) > $signed(cfar_cfar_cfarCore_rightThr); // @[FixedPointTypeClass.scala 55:59]
  assign cfar_cfar_cfarCore_greatestOf = cfar_cfar_cfarCore__T_70 ? $signed(cfar_cfar_cfarCore_leftThr) : $signed(cfar_cfar_cfarCore_rightThr); // @[CFARCoreWithMem.scala 143:23]
  assign cfar_cfar_cfarCore__T_71 = $signed(cfar_cfar_cfarCore_leftThr) < $signed(cfar_cfar_cfarCore_rightThr); // @[FixedPointTypeClass.scala 53:59]
  assign cfar_cfar_cfarCore_smallestOf = cfar_cfar_cfarCore__T_71 ? $signed(cfar_cfar_cfarCore_leftThr) : $signed(cfar_cfar_cfarCore_rightThr); // @[CFARCoreWithMem.scala 144:23]
  assign cfar_cfar_cfarCore__T_74 = $signed(cfar_cfar_cfarCore_rightThr) + $signed(cfar_cfar_cfarCore_leftThr); // @[FixedPointTypeClass.scala 20:58]
  assign cfar_cfar_cfarCore__T_75 = cfar_cfar_cfarCore__T_74[19:1]; // @[FixedPointTypeClass.scala 117:50]
  assign cfar_cfar_cfarCore__T_78 = 2'h1 == cfar_cfar_cfarCore_io_cfarMode; // @[Mux.scala 68:19]
  assign cfar_cfar_cfarCore__T_79 = cfar_cfar_cfarCore__T_78 ? $signed(cfar_cfar_cfarCore_greatestOf) : $signed(cfar_cfar_cfarCore_smallestOf); // @[Mux.scala 68:16]
  assign cfar_cfar_cfarCore__T_80 = 2'h0 == cfar_cfar_cfarCore_io_cfarMode; // @[Mux.scala 68:19]
  assign cfar_cfar_cfarCore_thrByModes = cfar_cfar_cfarCore__T_80 ? $signed({{1{cfar_cfar_cfarCore__T_75[18]}},cfar_cfar_cfarCore__T_75}) : $signed(cfar_cfar_cfarCore__T_79); // @[Mux.scala 68:16]
  assign cfar_cfar_cfarCore__T_81 = ~cfar_cfar_cfarCore_laggWindow_io_memFull; // @[CFARCoreWithMem.scala 152:9]
  assign cfar_cfar_cfarCore__T_83 = cfar_cfar_cfarCore__T_81 & cfar_cfar_cfarCore__T_47; // @[CFARCoreWithMem.scala 152:34]
  assign cfar_cfar_cfarCore__GEN_21 = cfar_cfar_cfarCore__T_83 | cfar_cfar_cfarCore_enableRightThr; // @[CFARCoreWithMem.scala 152:63]
  assign cfar_cfar_cfarCore__T_84 = ~cfar_cfar_cfarCore_leadWindow_io_memFull; // @[CFARCoreWithMem.scala 172:33]
  assign cfar_cfar_cfarCore__T_86 = cfar_cfar_cfarCore__T_84 & cfar_cfar_cfarCore__T_81; // @[CFARCoreWithMem.scala 172:56]
  assign cfar_cfar_cfarCore__T_90 = cfar_cfar_cfarCore_laggWindow_io_memFull & cfar_cfar_cfarCore__T_84; // @[CFARCoreWithMem.scala 174:57]
  assign cfar_cfar_cfarCore__T_91 = cfar_cfar_cfarCore_enableRightThr ? $signed(cfar_cfar_cfarCore_rightThr) : $signed(cfar_cfar_cfarCore_thrByModes); // @[CFARCoreWithMem.scala 177:36]
  assign cfar_cfar_cfarCore__T_92 = cfar_cfar_cfarCore__T_90 ? $signed(cfar_cfar_cfarCore_leftThr) : $signed(cfar_cfar_cfarCore__T_91); // @[CFARCoreWithMem.scala 174:34]
  assign cfar_cfar_cfarCore_thrWithoutScaling = cfar_cfar_cfarCore__T_86 ? $signed(20'sh0) : $signed(cfar_cfar_cfarCore__T_92); // @[CFARCoreWithMem.scala 172:32]
  assign cfar_cfar_cfarCore__GEN_51 = {{4{cfar_cfar_cfarCore_io_thresholdScaler[15]}},cfar_cfar_cfarCore_io_thresholdScaler}; // @[FixedPointTypeClass.scala 211:35]
  assign cfar_cfar_cfarCore_threshold = cfar_cfar_cfarCore__T_94[35:13]; // @[FixedPointTypeClass.scala 153:43]
  assign cfar_cfar_cfarCore__T_96 = cfar_cfar_cfarCore_io_guardCells - 4'h1; // @[CFARCoreWithMem.scala 197:74]
  assign cfar_cfar_cfarCore__T_97 = cfar_cfar_cfarCore__T_96[2:0];
  assign cfar_cfar_cfarCore__GEN_25 = cfar_cfar_cfarCore_laggGuard_io_parallelOut_0; // @[Reg.scala 16:23]
  assign cfar_cfar_cfarCore__T_98 = $signed(cfar_cfar_cfarCore_cutDelayed) > $signed(cfar_cfar_cfarCore_leftNeighb); // @[FixedPointTypeClass.scala 55:59]
  assign cfar_cfar_cfarCore__T_99 = $signed(cfar_cfar_cfarCore_cutDelayed) > $signed(cfar_cfar_cfarCore_rightNeighb); // @[FixedPointTypeClass.scala 55:59]
  assign cfar_cfar_cfarCore_isLocalMax = cfar_cfar_cfarCore__T_98 & cfar_cfar_cfarCore__T_99; // @[CFARCoreWithMem.scala 199:44]
  assign cfar_cfar_cfarCore__GEN_52 = {$signed(cfar_cfar_cfarCore_cutDelayed), 1'h0}; // @[FixedPointTypeClass.scala 55:59]
  assign cfar_cfar_cfarCore__GEN_53 = {{6{cfar_cfar_cfarCore__GEN_52[16]}},cfar_cfar_cfarCore__GEN_52}; // @[FixedPointTypeClass.scala 55:59]
  assign cfar_cfar_cfarCore_isPeak = $signed(cfar_cfar_cfarCore__GEN_53) > $signed(cfar_cfar_cfarCore_threshold); // @[FixedPointTypeClass.scala 55:59]
  assign cfar_cfar_cfarCore__T_100 = ~cfar_cfar_cfarCore_initialInDone; // @[CFARCoreWithMem.scala 216:20]
  assign cfar_cfar_cfarCore__T_101 = ~cfar_cfar_cfarCore_flushingDelayed; // @[CFARCoreWithMem.scala 216:54]
  assign cfar_cfar_cfarCore__T_102 = cfar_cfar_cfarCore_io_out_ready & cfar_cfar_cfarCore__T_101; // @[CFARCoreWithMem.scala 216:51]
  assign cfar_cfar_cfarCore__T_108 = cfar_cfar_cfarCore_flushingDelayed & cfar_cfar_cfarCore__T_107; // @[CFARCoreWithMem.scala 218:123]
  assign cfar_cfar_cfarCore__T_110 = cfar_cfar_cfarCore_isPeak & cfar_cfar_cfarCore_isLocalMax; // @[CFARCoreWithMem.scala 223:63]
  assign cfar_cfar_cfarCore__T_122 = cfar_cfar_cfarCore_flushingDelayed & cfar_cfar_cfarCore__T_121; // @[CFARCoreWithMem.scala 231:123]
  assign cfar_cfar_cfarCore_io_in_ready = cfar_cfar_cfarCore__T_100 | cfar_cfar_cfarCore__T_102; // @[CFARCoreWithMem.scala 41:20 CFARCoreWithMem.scala 216:17]
  assign cfar_cfar_cfarCore_io_out_valid = cfar_cfar_cfarCore_Queue_io_deq_valid; // @[CFARCoreWithMem.scala 241:18]
  assign cfar_cfar_cfarCore_io_out_bits_peak = cfar_cfar_cfarCore_Queue_io_deq_bits_peak; // @[CFARCoreWithMem.scala 239:22]
  assign cfar_cfar_cfarCore_io_out_bits_cut = cfar_cfar_cfarCore_Queue_io_deq_bits_cut; // @[CFARCoreWithMem.scala 238:27]
  assign cfar_cfar_cfarCore_io_out_bits_threshold = cfar_cfar_cfarCore_Queue_io_deq_bits_threshold; // @[CFARCoreWithMem.scala 240:27]
  assign cfar_cfar_cfarCore_io_lastOut = cfar_cfar_cfarCore_Queue_2_io_deq_bits; // @[CFARCoreWithMem.scala 235:16]
  assign cfar_cfar_cfarCore_io_fftBin = cfar_cfar_cfarCore_cntOut; // @[CFARCoreWithMem.scala 242:15]
  assign cfar_cfar_cfarCore_laggWindow_clock = cfar_cfar_cfarCore_clock;
  assign cfar_cfar_cfarCore_laggWindow_reset = cfar_cfar_cfarCore_reset;
  assign cfar_cfar_cfarCore_laggWindow_io_depth = cfar_cfar_cfarCore_io_windowCells; // @[CFARCoreWithMem.scala 42:23]
  assign cfar_cfar_cfarCore_laggWindow_io_in_valid = cfar_cfar_cfarCore_io_in_valid; // @[CFARCoreWithMem.scala 41:20]
  assign cfar_cfar_cfarCore_laggWindow_io_in_bits = cfar_cfar_cfarCore_io_in_bits; // @[CFARCoreWithMem.scala 41:20]
  assign cfar_cfar_cfarCore_laggWindow_io_lastIn = cfar_cfar_cfarCore_io_lastIn; // @[CFARCoreWithMem.scala 43:24]
  assign cfar_cfar_cfarCore_laggWindow_io_out_ready = cfar_cfar_cfarCore_laggGuard_io_in_ready; // @[CFARCoreWithMem.scala 46:19]
  assign cfar_cfar_cfarCore_laggGuard_clock = cfar_cfar_cfarCore_clock;
  assign cfar_cfar_cfarCore_laggGuard_reset = cfar_cfar_cfarCore_reset;
  assign cfar_cfar_cfarCore_laggGuard_io_depth = cfar_cfar_cfarCore_io_guardCells; // @[CFARCoreWithMem.scala 48:23]
  assign cfar_cfar_cfarCore_laggGuard_io_in_valid = cfar_cfar_cfarCore_laggWindow_io_out_valid; // @[CFARCoreWithMem.scala 46:19]
  assign cfar_cfar_cfarCore_laggGuard_io_in_bits = cfar_cfar_cfarCore_laggWindow_io_out_bits; // @[CFARCoreWithMem.scala 46:19]
  assign cfar_cfar_cfarCore_laggGuard_io_lastIn = cfar_cfar_cfarCore_laggWindow_io_lastOut; // @[CFARCoreWithMem.scala 47:23]
  assign cfar_cfar_cfarCore_laggGuard_io_out_ready = cfar_cfar_cfarCore_cellUnderTest_io_in_ready; // @[CFARCoreWithMem.scala 51:23]
  assign cfar_cfar_cfarCore_cellUnderTest_clock = cfar_cfar_cfarCore_clock;
  assign cfar_cfar_cfarCore_cellUnderTest_reset = cfar_cfar_cfarCore_reset;
  assign cfar_cfar_cfarCore_cellUnderTest_io_in_valid = cfar_cfar_cfarCore_laggGuard_io_out_valid; // @[CFARCoreWithMem.scala 51:23]
  assign cfar_cfar_cfarCore_cellUnderTest_io_in_bits = cfar_cfar_cfarCore_laggGuard_io_out_bits; // @[CFARCoreWithMem.scala 51:23]
  assign cfar_cfar_cfarCore_cellUnderTest_io_lastIn = cfar_cfar_cfarCore_laggGuard_io_lastOut; // @[CFARCoreWithMem.scala 52:27]
  assign cfar_cfar_cfarCore_cellUnderTest_io_out_ready = cfar_cfar_cfarCore_leadWindow_io_memFull ? cfar_cfar_cfarCore_leadWindow_io_in_ready : cfar_cfar_cfarCore_io_out_ready; // @[CFARCoreWithMem.scala 56:19 CFARCoreWithMem.scala 71:30]
  assign cfar_cfar_cfarCore_leadGuard_clock = cfar_cfar_cfarCore_clock;
  assign cfar_cfar_cfarCore_leadGuard_reset = cfar_cfar_cfarCore_reset;
  assign cfar_cfar_cfarCore_leadGuard_io_depth = cfar_cfar_cfarCore_io_guardCells; // @[CFARCoreWithMem.scala 57:22]
  assign cfar_cfar_cfarCore_leadGuard_io_in_valid = cfar_cfar_cfarCore_cellUnderTest_io_out_valid; // @[CFARCoreWithMem.scala 56:19]
  assign cfar_cfar_cfarCore_leadGuard_io_in_bits = cfar_cfar_cfarCore_cellUnderTest_io_out_bits; // @[CFARCoreWithMem.scala 56:19]
  assign cfar_cfar_cfarCore_leadGuard_io_lastIn = cfar_cfar_cfarCore_cellUnderTest_io_lastOut; // @[CFARCoreWithMem.scala 58:23]
  assign cfar_cfar_cfarCore_leadGuard_io_out_ready = cfar_cfar_cfarCore_leadWindow_io_in_ready; // @[CFARCoreWithMem.scala 61:26 CFARCoreWithMem.scala 65:20]
  assign cfar_cfar_cfarCore_leadWindow_clock = cfar_cfar_cfarCore_clock;
  assign cfar_cfar_cfarCore_leadWindow_reset = cfar_cfar_cfarCore_reset;
  assign cfar_cfar_cfarCore_leadWindow_io_depth = cfar_cfar_cfarCore_io_windowCells; // @[CFARCoreWithMem.scala 64:23]
  assign cfar_cfar_cfarCore_leadWindow_io_in_valid = cfar_cfar_cfarCore_leadGuard_io_out_valid; // @[CFARCoreWithMem.scala 65:20]
  assign cfar_cfar_cfarCore_leadWindow_io_in_bits = cfar_cfar_cfarCore_leadGuard_io_out_bits; // @[CFARCoreWithMem.scala 65:20]
  assign cfar_cfar_cfarCore_leadWindow_io_lastIn = cfar_cfar_cfarCore_leadGuard_io_lastOut; // @[CFARCoreWithMem.scala 72:24]
  assign cfar_cfar_cfarCore_leadWindow_io_out_ready = cfar_cfar_cfarCore_io_out_ready; // @[CFARCoreWithMem.scala 69:27]
  assign cfar_cfar_cfarCore_Queue_clock = cfar_cfar_cfarCore_clock;
  assign cfar_cfar_cfarCore_Queue_reset = cfar_cfar_cfarCore_reset;
  assign cfar_cfar_cfarCore_Queue_io_enq_valid = cfar_cfar_cfarCore__T_106 | cfar_cfar_cfarCore__T_108; // @[CFARCoreWithMem.scala 218:28]
  assign cfar_cfar_cfarCore_Queue_io_enq_bits_peak = cfar_cfar_cfarCore_io_peakGrouping ? cfar_cfar_cfarCore__T_110 : cfar_cfar_cfarCore_isPeak; // @[CFARCoreWithMem.scala 223:32]
  assign cfar_cfar_cfarCore_Queue_io_enq_bits_cut = cfar_cfar_cfarCore_cutDelayed; // @[CFARCoreWithMem.scala 221:37]
  assign cfar_cfar_cfarCore__GEN_55 = cfar_cfar_cfarCore_threshold[22:1]; // @[CFARCoreWithMem.scala 222:37]
  assign cfar_cfar_cfarCore_Queue_io_enq_bits_threshold = cfar_cfar_cfarCore__GEN_55[15:0]; // @[CFARCoreWithMem.scala 222:37]
  assign cfar_cfar_cfarCore_Queue_io_deq_ready = cfar_cfar_cfarCore_io_out_ready; // @[CFARCoreWithMem.scala 224:28]
  assign cfar_cfar_cfarCore_Queue_2_clock = cfar_cfar_cfarCore_clock;
  assign cfar_cfar_cfarCore_Queue_2_reset = cfar_cfar_cfarCore_reset;
  assign cfar_cfar_cfarCore_Queue_2_io_enq_valid = cfar_cfar_cfarCore__T_120 | cfar_cfar_cfarCore__T_122; // @[CFARCoreWithMem.scala 231:28]
  assign cfar_cfar_cfarCore_Queue_2_io_enq_bits = cfar_cfar_cfarCore_lastOut; // @[CFARCoreWithMem.scala 232:27]
  assign cfar_cfar_cfarCore_Queue_2_io_deq_ready = cfar_cfar_cfarCore_io_out_ready; // @[CFARCoreWithMem.scala 234:28]
  assign cfar_cfar_io_in_ready = cfar_cfar_cfarCore_io_in_ready; // @[CFARcore.scala 68:18]
  assign cfar_cfar_io_out_valid = cfar_cfar_cfarCore_io_out_valid; // @[CFARcore.scala 95:19]
  assign cfar_cfar_io_out_bits_peak = cfar_cfar_cfarCore_io_out_bits_peak; // @[CFARcore.scala 95:19]
  assign cfar_cfar_io_out_bits_cut = cfar_cfar_cfarCore_io_out_bits_cut; // @[CFARcore.scala 95:19]
  assign cfar_cfar_io_out_bits_threshold = cfar_cfar_cfarCore_io_out_bits_threshold; // @[CFARcore.scala 95:19]
  assign cfar_cfar_io_lastOut = cfar_cfar_cfarCore_io_lastOut; // @[CFARcore.scala 96:14]
  assign cfar_cfar_io_fftBin = cfar_cfar_cfarCore_io_fftBin; // @[CFARcore.scala 97:13]
  assign cfar_cfar_cfarCore_clock = cfar_cfar_clock;
  assign cfar_cfar_cfarCore_reset = cfar_cfar_reset;
  assign cfar_cfar_cfarCore_io_in_valid = cfar_cfar_io_in_valid; // @[CFARcore.scala 68:18]
  assign cfar_cfar_cfarCore_io_in_bits = cfar_cfar_io_in_bits; // @[CFARcore.scala 68:18]
  assign cfar_cfar_cfarCore_io_lastIn = cfar_cfar_io_lastIn; // @[CFARcore.scala 69:22]
  assign cfar_cfar_cfarCore_io_fftWin = cfar_cfar_io_fftWin; // @[CFARcore.scala 70:22]
  assign cfar_cfar_cfarCore_io_thresholdScaler = cfar_cfar_io_thresholdScaler; // @[CFARcore.scala 71:31]
  assign cfar_cfar_cfarCore_io_divSum = cfar_cfar_io_divSum; // @[CFARcore.scala 77:28]
  assign cfar_cfar_cfarCore_io_peakGrouping = cfar_cfar_io_peakGrouping; // @[CFARcore.scala 79:28]
  assign cfar_cfar_cfarCore_io_cfarMode = cfar_cfar_io_cfarMode; // @[CFARcore.scala 83:24]
  assign cfar_cfar_cfarCore_io_windowCells = cfar_cfar_io_windowCells; // @[CFARcore.scala 84:27]
  assign cfar_cfar_cfarCore_io_guardCells = cfar_cfar_io_guardCells; // @[CFARcore.scala 85:26]
  assign cfar_cfar_cfarCore_io_out_ready = cfar_cfar_io_out_ready; // @[CFARcore.scala 95:19]
  assign cfar_Queue__T_read__T_18_addr = cfar_Queue_value_1;
  assign cfar_Queue__T_read__T_18_data = cfar_Queue__T_read[cfar_Queue__T_read__T_18_addr]; // @[Decoupled.scala 209:24]
  assign cfar_Queue__T_read__T_10_data = cfar_Queue_io_enq_bits_read;
  assign cfar_Queue__T_read__T_10_addr = cfar_Queue_value;
  assign cfar_Queue__T_read__T_10_mask = 1'h1;
  assign cfar_Queue__T_read__T_10_en = cfar_Queue_io_enq_ready & cfar_Queue_io_enq_valid;
  assign cfar_Queue__T_data__T_18_addr = cfar_Queue_value_1;
  assign cfar_Queue__T_data__T_18_data = cfar_Queue__T_data[cfar_Queue__T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign cfar_Queue__T_data__T_10_data = cfar_Queue_io_enq_bits_data;
  assign cfar_Queue__T_data__T_10_addr = cfar_Queue_value;
  assign cfar_Queue__T_data__T_10_mask = 1'h1;
  assign cfar_Queue__T_data__T_10_en = cfar_Queue_io_enq_ready & cfar_Queue_io_enq_valid;
  assign cfar_Queue__T_extra__T_18_addr = cfar_Queue_value_1;
  assign cfar_Queue__T_extra__T_18_data = cfar_Queue__T_extra[cfar_Queue__T_extra__T_18_addr]; // @[Decoupled.scala 209:24]
  assign cfar_Queue__T_extra__T_10_data = cfar_Queue_io_enq_bits_extra;
  assign cfar_Queue__T_extra__T_10_addr = cfar_Queue_value;
  assign cfar_Queue__T_extra__T_10_mask = 1'h1;
  assign cfar_Queue__T_extra__T_10_en = cfar_Queue_io_enq_ready & cfar_Queue_io_enq_valid;
  assign cfar_Queue__T_2 = cfar_Queue_value == cfar_Queue_value_1; // @[Decoupled.scala 214:41]
  assign cfar_Queue__T_3 = ~cfar_Queue__T_1; // @[Decoupled.scala 215:36]
  assign cfar_Queue__T_4 = cfar_Queue__T_2 & cfar_Queue__T_3; // @[Decoupled.scala 215:33]
  assign cfar_Queue__T_5 = cfar_Queue__T_2 & cfar_Queue__T_1; // @[Decoupled.scala 216:32]
  assign cfar_Queue__T_6 = cfar_Queue_io_enq_ready & cfar_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign cfar_Queue__T_8 = cfar_Queue_io_deq_ready & cfar_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign cfar_Queue__T_12 = cfar_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign cfar_Queue__T_14 = cfar_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign cfar_Queue__T_15 = cfar_Queue__T_6 != cfar_Queue__T_8; // @[Decoupled.scala 227:16]
  assign cfar_Queue_io_enq_ready = ~cfar_Queue__T_5; // @[Decoupled.scala 232:16]
  assign cfar_Queue_io_deq_valid = ~cfar_Queue__T_4; // @[Decoupled.scala 231:16]
  assign cfar_Queue_io_deq_bits_read = cfar_Queue__T_read__T_18_data; // @[Decoupled.scala 233:15]
  assign cfar_Queue_io_deq_bits_data = cfar_Queue__T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign cfar_Queue_io_deq_bits_extra = cfar_Queue__T_extra__T_18_data; // @[Decoupled.scala 233:15]
  assign cfar__T_11 = {cfar_cfar_io_out_bits_threshold,cfar_cfar_io_out_bits_cut,cfar_cfar_io_fftBin,cfar_cfar_io_out_bits_peak}; // @[Cat.scala 29:58]
  assign cfar__T_13 = cfar_auto_mem_in_aw_valid & cfar_auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign cfar__T_14 = cfar_auto_mem_in_ar_valid | cfar__T_13; // @[RegisterRouter.scala 40:26]
  assign cfar__T_15 = ~cfar_auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign cfar__T_58_ready = cfar_Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign cfar__T_22 = cfar_auto_mem_in_ar_valid ? cfar_auto_mem_in_ar_bits_addr : cfar_auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign cfar__T_56 = cfar__T_22[29:2]; // @[RegisterRouter.scala 52:27]
  assign cfar__T_12_bits_index = cfar__T_56[5:0]; // @[RegisterRouter.scala 37:18 RegisterRouter.scala 52:19]
  assign cfar__T_282 = cfar__T_12_bits_index[2]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_281 = cfar__T_12_bits_index[1]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_280 = cfar__T_12_bits_index[0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_287 = {cfar__T_282,cfar__T_281,cfar__T_280}; // @[Cat.scala 29:58]
  assign cfar__T_62 = cfar__T_12_bits_index & 6'h38; // @[RegisterRouter.scala 59:16]
  assign cfar__T_70 = cfar__T_62 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign cfar__T_16 = cfar__T_58_ready & cfar__T_15; // @[RegisterRouter.scala 42:26]
  assign cfar__T_24 = cfar_auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 64:49]
  assign cfar__T_25 = 2'h1 << cfar__T_24; // @[OneHot.scala 65:12]
  assign cfar__T_27 = cfar__T_25 | 2'h1; // @[Misc.scala 200:81]
  assign cfar__T_28 = cfar_auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign cfar__T_29 = cfar__T_27[1]; // @[Misc.scala 207:26]
  assign cfar__T_30 = cfar_auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 208:26]
  assign cfar__T_31 = ~cfar__T_30; // @[Misc.scala 209:20]
  assign cfar__T_33 = cfar__T_29 & cfar__T_31; // @[Misc.scala 213:38]
  assign cfar__T_34 = cfar__T_28 | cfar__T_33; // @[Misc.scala 213:29]
  assign cfar__T_36 = cfar__T_29 & cfar__T_30; // @[Misc.scala 213:38]
  assign cfar__T_37 = cfar__T_28 | cfar__T_36; // @[Misc.scala 213:29]
  assign cfar__T_38 = cfar__T_27[0]; // @[Misc.scala 207:26]
  assign cfar__T_39 = cfar_auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 208:26]
  assign cfar__T_40 = ~cfar__T_39; // @[Misc.scala 209:20]
  assign cfar__T_41 = cfar__T_31 & cfar__T_40; // @[Misc.scala 212:27]
  assign cfar__T_42 = cfar__T_38 & cfar__T_41; // @[Misc.scala 213:38]
  assign cfar__T_43 = cfar__T_34 | cfar__T_42; // @[Misc.scala 213:29]
  assign cfar__T_44 = cfar__T_31 & cfar__T_39; // @[Misc.scala 212:27]
  assign cfar__T_45 = cfar__T_38 & cfar__T_44; // @[Misc.scala 213:38]
  assign cfar__T_46 = cfar__T_34 | cfar__T_45; // @[Misc.scala 213:29]
  assign cfar__T_47 = cfar__T_30 & cfar__T_40; // @[Misc.scala 212:27]
  assign cfar__T_48 = cfar__T_38 & cfar__T_47; // @[Misc.scala 213:38]
  assign cfar__T_49 = cfar__T_37 | cfar__T_48; // @[Misc.scala 213:29]
  assign cfar__T_50 = cfar__T_30 & cfar__T_39; // @[Misc.scala 212:27]
  assign cfar__T_51 = cfar__T_38 & cfar__T_50; // @[Misc.scala 213:38]
  assign cfar__T_52 = cfar__T_37 | cfar__T_51; // @[Misc.scala 213:29]
  assign cfar__T_55 = {cfar__T_52,cfar__T_49,cfar__T_46,cfar__T_43}; // @[Cat.scala 29:58]
  assign cfar__T_57 = cfar_auto_mem_in_ar_valid ? cfar__T_55 : cfar_auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign cfar__T_81 = cfar__T_57[0]; // @[Bitwise.scala 26:51]
  assign cfar__T_82 = cfar__T_57[1]; // @[Bitwise.scala 26:51]
  assign cfar__T_83 = cfar__T_57[2]; // @[Bitwise.scala 26:51]
  assign cfar__T_84 = cfar__T_57[3]; // @[Bitwise.scala 26:51]
  assign cfar__T_86 = cfar__T_81 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign cfar__T_88 = cfar__T_82 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign cfar__T_90 = cfar__T_83 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign cfar__T_92 = cfar__T_84 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign cfar__T_95 = {cfar__T_92,cfar__T_90,cfar__T_88,cfar__T_86}; // @[Cat.scala 29:58]
  assign cfar__T_111 = cfar__T_95[9:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_114 = cfar__T_111 == 10'h3ff; // @[RegisterRouter.scala 59:16]
  assign cfar__T_306 = cfar__T_14 & cfar__T_58_ready; // @[RegisterRouter.scala 59:16]
  assign cfar__T_288 = 8'h1 << cfar__T_287; // @[OneHot.scala 58:35]
  assign cfar__T_289 = cfar__T_288[0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_353 = cfar__T_306 & cfar__T_15; // @[RegisterRouter.scala 59:16]
  assign cfar__T_355 = cfar__T_353 & cfar__T_289; // @[RegisterRouter.scala 59:16]
  assign cfar__T_356 = cfar__T_355 & cfar__T_70; // @[RegisterRouter.scala 59:16]
  assign cfar__T_121 = cfar__T_356 & cfar__T_114; // @[RegisterRouter.scala 59:16]
  assign cfar__T_123 = cfar_auto_mem_in_w_bits_data[9:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_134 = cfar__T_95[3:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_137 = cfar__T_134 == 4'hf; // @[RegisterRouter.scala 59:16]
  assign cfar__T_294 = cfar__T_288[5]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_380 = cfar__T_353 & cfar__T_294; // @[RegisterRouter.scala 59:16]
  assign cfar__T_381 = cfar__T_380 & cfar__T_70; // @[RegisterRouter.scala 59:16]
  assign cfar__T_144 = cfar__T_381 & cfar__T_137; // @[RegisterRouter.scala 59:16]
  assign cfar__T_146 = cfar_auto_mem_in_w_bits_data[3:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_157 = cfar__T_95[15:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_160 = cfar__T_157 == 16'hffff; // @[RegisterRouter.scala 59:16]
  assign cfar__T_290 = cfar__T_288[1]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_360 = cfar__T_353 & cfar__T_290; // @[RegisterRouter.scala 59:16]
  assign cfar__T_361 = cfar__T_360 & cfar__T_70; // @[RegisterRouter.scala 59:16]
  assign cfar__T_167 = cfar__T_361 & cfar__T_160; // @[RegisterRouter.scala 59:16]
  assign cfar__T_169 = cfar_auto_mem_in_w_bits_data[15:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_180 = cfar__T_95[2:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_183 = cfar__T_180 == 3'h7; // @[RegisterRouter.scala 59:16]
  assign cfar__T_295 = cfar__T_288[6]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_385 = cfar__T_353 & cfar__T_295; // @[RegisterRouter.scala 59:16]
  assign cfar__T_386 = cfar__T_385 & cfar__T_70; // @[RegisterRouter.scala 59:16]
  assign cfar__T_190 = cfar__T_386 & cfar__T_183; // @[RegisterRouter.scala 59:16]
  assign cfar__T_192 = cfar_auto_mem_in_w_bits_data[2:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_203 = cfar__T_95[0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_291 = cfar__T_288[2]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_365 = cfar__T_353 & cfar__T_291; // @[RegisterRouter.scala 59:16]
  assign cfar__T_366 = cfar__T_365 & cfar__T_70; // @[RegisterRouter.scala 59:16]
  assign cfar__T_213 = cfar__T_366 & cfar__T_203; // @[RegisterRouter.scala 59:16]
  assign cfar__T_215 = cfar_auto_mem_in_w_bits_data[0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_226 = cfar__T_95[1:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_229 = cfar__T_226 == 2'h3; // @[RegisterRouter.scala 59:16]
  assign cfar__T_292 = cfar__T_288[3]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_370 = cfar__T_353 & cfar__T_292; // @[RegisterRouter.scala 59:16]
  assign cfar__T_371 = cfar__T_370 & cfar__T_70; // @[RegisterRouter.scala 59:16]
  assign cfar__T_236 = cfar__T_371 & cfar__T_229; // @[RegisterRouter.scala 59:16]
  assign cfar__T_238 = cfar_auto_mem_in_w_bits_data[1:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_249 = cfar__T_95[6:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_252 = cfar__T_249 == 7'h7f; // @[RegisterRouter.scala 59:16]
  assign cfar__T_293 = cfar__T_288[4]; // @[RegisterRouter.scala 59:16]
  assign cfar__T_375 = cfar__T_353 & cfar__T_293; // @[RegisterRouter.scala 59:16]
  assign cfar__T_376 = cfar__T_375 & cfar__T_70; // @[RegisterRouter.scala 59:16]
  assign cfar__T_259 = cfar__T_376 & cfar__T_252; // @[RegisterRouter.scala 59:16]
  assign cfar__T_261 = cfar_auto_mem_in_w_bits_data[6:0]; // @[RegisterRouter.scala 59:16]
  assign cfar__GEN_40 = 3'h1 == cfar__T_287 ? cfar__T_70 : cfar__T_70; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_41 = 3'h2 == cfar__T_287 ? cfar__T_70 : cfar__GEN_40; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_42 = 3'h3 == cfar__T_287 ? cfar__T_70 : cfar__GEN_41; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_43 = 3'h4 == cfar__T_287 ? cfar__T_70 : cfar__GEN_42; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_44 = 3'h5 == cfar__T_287 ? cfar__T_70 : cfar__GEN_43; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_45 = 3'h6 == cfar__T_287 ? cfar__T_70 : cfar__GEN_44; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_55 = 3'h7 == cfar__T_287; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_46 = cfar__GEN_55 | cfar__GEN_45; // @[MuxLiteral.scala 48:10]
  assign cfar__T_498_0 = {{6'd0}, cfar_fftWin}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign cfar__GEN_48 = 3'h1 == cfar__T_287 ? cfar_thresholdScaler : cfar__T_498_0; // @[MuxLiteral.scala 48:10]
  assign cfar__T_498_2 = {{15'd0}, cfar_peakGrouping}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign cfar__GEN_49 = 3'h2 == cfar__T_287 ? cfar__T_498_2 : cfar__GEN_48; // @[MuxLiteral.scala 48:10]
  assign cfar__T_498_3 = {{14'd0}, cfar_cfarMode}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign cfar__GEN_50 = 3'h3 == cfar__T_287 ? cfar__T_498_3 : cfar__GEN_49; // @[MuxLiteral.scala 48:10]
  assign cfar__T_498_4 = {{9'd0}, cfar_windowCells}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign cfar__GEN_51 = 3'h4 == cfar__T_287 ? cfar__T_498_4 : cfar__GEN_50; // @[MuxLiteral.scala 48:10]
  assign cfar__T_498_5 = {{12'd0}, cfar_guardCells}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign cfar__GEN_52 = 3'h5 == cfar__T_287 ? cfar__T_498_5 : cfar__GEN_51; // @[MuxLiteral.scala 48:10]
  assign cfar__T_498_6 = {{13'd0}, cfar__T_6}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign cfar__GEN_53 = 3'h6 == cfar__T_287 ? cfar__T_498_6 : cfar__GEN_52; // @[MuxLiteral.scala 48:10]
  assign cfar__GEN_54 = 3'h7 == cfar__T_287 ? 16'h0 : cfar__GEN_53; // @[MuxLiteral.scala 48:10]
  assign cfar__T_500 = cfar__GEN_46 ? cfar__GEN_54 : 16'h0; // @[RegisterRouter.scala 59:16]
  assign cfar__T_501_bits_read = cfar_Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign cfar__T_501_valid = cfar_Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign cfar__T_504 = ~cfar__T_501_bits_read; // @[RegisterRouter.scala 65:29]
  assign cfar_auto_mem_in_aw_ready = cfar__T_16 & cfar_auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign cfar_auto_mem_in_w_ready = cfar__T_16 & cfar_auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign cfar_auto_mem_in_b_valid = cfar__T_501_valid & cfar__T_504; // @[LazyModule.scala 173:31]
  assign cfar_auto_mem_in_b_bits_id = cfar_Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign cfar_auto_mem_in_ar_ready = cfar_Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign cfar_auto_mem_in_r_valid = cfar__T_501_valid & cfar__T_501_bits_read; // @[LazyModule.scala 173:31]
  assign cfar_auto_mem_in_r_bits_id = cfar_Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign cfar_auto_mem_in_r_bits_data = cfar_Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign cfar_auto_master_out_valid = cfar_cfar_io_out_valid; // @[LazyModule.scala 173:49]
  assign cfar_auto_master_out_bits_data = {{6'd0}, cfar__T_11}; // @[LazyModule.scala 173:49]
  assign cfar_auto_master_out_bits_last = cfar_cfar_io_lastOut; // @[LazyModule.scala 173:49]
  assign cfar_auto_slave_in_ready = cfar_cfar_io_in_ready; // @[LazyModule.scala 173:31]
  assign cfar_cfar_clock = cfar_clock;
  assign cfar_cfar_reset = cfar_reset;
  assign cfar_cfar_io_in_valid = cfar_auto_slave_in_valid; // @[CFARDspBlock.scala 97:22]
  assign cfar_cfar_io_in_bits = cfar_auto_slave_in_bits_data; // @[CFARDspBlock.scala 98:21]
  assign cfar_cfar_io_lastIn = cfar_auto_slave_in_bits_last; // @[CFARDspBlock.scala 135:25]
  assign cfar_cfar_io_fftWin = cfar_fftWin; // @[CFARDspBlock.scala 100:20]
  assign cfar_cfar_io_thresholdScaler = cfar_thresholdScaler; // @[CFARDspBlock.scala 101:29]
  assign cfar_cfar_io_divSum = cfar__T_6; // @[CFARDspBlock.scala 112:26]
  assign cfar_cfar_io_peakGrouping = cfar_peakGrouping; // @[CFARDspBlock.scala 124:26]
  assign cfar_cfar_io_cfarMode = cfar_cfarMode; // @[CFARDspBlock.scala 132:25]
  assign cfar_cfar_io_windowCells = cfar_windowCells; // @[CFARDspBlock.scala 133:25]
  assign cfar_cfar_io_guardCells = cfar_guardCells; // @[CFARDspBlock.scala 134:25]
  assign cfar_cfar_io_out_ready = cfar_auto_master_out_ready; // @[CFARDspBlock.scala 162:24]
  assign cfar_Queue_clock = cfar_clock;
  assign cfar_Queue_reset = cfar_reset;
  assign cfar_Queue_io_enq_valid = cfar_auto_mem_in_ar_valid | cfar__T_13; // @[Decoupled.scala 288:22]
  assign cfar_Queue_io_enq_bits_read = cfar_auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign cfar_Queue_io_enq_bits_data = {{16'd0}, cfar__T_500}; // @[Decoupled.scala 289:21]
  assign cfar_Queue_io_enq_bits_extra = cfar_auto_mem_in_ar_valid ? cfar_auto_mem_in_ar_bits_id : cfar_auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign cfar_Queue_io_deq_ready = cfar__T_501_bits_read ? cfar_auto_mem_in_r_ready : cfar_auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
  assign widthAdapter_1__T = widthAdapter_1_auto_in_bits_data[15:0]; // @[AXI4StreamWidthAdapter.scala 154:10]
  assign widthAdapter_1__T_1 = widthAdapter_1_auto_in_bits_data[31:16]; // @[AXI4StreamWidthAdapter.scala 154:10]
  assign widthAdapter_1__T_2 = widthAdapter_1_auto_in_bits_data[47:32]; // @[AXI4StreamWidthAdapter.scala 154:10]
  assign widthAdapter_1__T_5 = widthAdapter_1_auto_in_valid & widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 159:14]
  assign widthAdapter_1__T_6 = widthAdapter_1__T_4 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign widthAdapter_1__T_7 = widthAdapter_1__T_4 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign widthAdapter_1__T_8 = widthAdapter_1__T_6 ? 3'h0 : widthAdapter_1__T_7; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign widthAdapter_1__GEN_0 = widthAdapter_1__T_5 ? widthAdapter_1__T_8 : {{1'd0}, widthAdapter_1__T_4}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign widthAdapter_1_ir0 = widthAdapter_1__T_6 & widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign widthAdapter_1__T_12 = widthAdapter_1__T_10 == 2'h2; // @[AXI4StreamWidthAdapter.scala 168:38]
  assign widthAdapter_1__T_13 = widthAdapter_1__T_10 + 2'h1; // @[AXI4StreamWidthAdapter.scala 168:60]
  assign widthAdapter_1__T_14 = widthAdapter_1__T_12 ? 3'h0 : widthAdapter_1__T_13; // @[AXI4StreamWidthAdapter.scala 168:33]
  assign widthAdapter_1__GEN_1 = widthAdapter_1__T_5 ? widthAdapter_1__T_14 : {{1'd0}, widthAdapter_1__T_10}; // @[AXI4StreamWidthAdapter.scala 168:21]
  assign widthAdapter_1_ir1 = widthAdapter_1__T_12 & widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 170:60]
  assign widthAdapter_1__T_21 = widthAdapter_1__T_19 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign widthAdapter_1__T_22 = widthAdapter_1__T_19 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign widthAdapter_1__T_23 = widthAdapter_1__T_21 ? 3'h0 : widthAdapter_1__T_22; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign widthAdapter_1__GEN_2 = widthAdapter_1__T_5 ? widthAdapter_1__T_23 : {{1'd0}, widthAdapter_1__T_19}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign widthAdapter_1_ir2 = widthAdapter_1__T_21 & widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign widthAdapter_1__T_28 = widthAdapter_1__T_26 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign widthAdapter_1__T_29 = widthAdapter_1__T_26 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign widthAdapter_1__T_30 = widthAdapter_1__T_28 ? 3'h0 : widthAdapter_1__T_29; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign widthAdapter_1__GEN_3 = widthAdapter_1__T_5 ? widthAdapter_1__T_30 : {{1'd0}, widthAdapter_1__T_26}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign widthAdapter_1_ir3 = widthAdapter_1__T_28 & widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign widthAdapter_1__T_35 = widthAdapter_1__T_33 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign widthAdapter_1__T_36 = widthAdapter_1__T_33 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign widthAdapter_1__T_37 = widthAdapter_1__T_35 ? 3'h0 : widthAdapter_1__T_36; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign widthAdapter_1__GEN_4 = widthAdapter_1__T_5 ? widthAdapter_1__T_37 : {{1'd0}, widthAdapter_1__T_33}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign widthAdapter_1_ir4 = widthAdapter_1__T_35 & widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign widthAdapter_1__T_55 = widthAdapter_1_ir0 == widthAdapter_1_ir1; // @[AXI4StreamWidthAdapter.scala 46:16]
  assign widthAdapter_1__T_57 = widthAdapter_1__T_55 | widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign widthAdapter_1__T_58 = ~widthAdapter_1__T_57; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign widthAdapter_1__T_59 = widthAdapter_1_ir0 == widthAdapter_1_ir2; // @[AXI4StreamWidthAdapter.scala 47:16]
  assign widthAdapter_1__T_61 = widthAdapter_1__T_59 | widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign widthAdapter_1__T_62 = ~widthAdapter_1__T_61; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign widthAdapter_1__T_63 = widthAdapter_1_ir0 == widthAdapter_1_ir3; // @[AXI4StreamWidthAdapter.scala 48:16]
  assign widthAdapter_1__T_65 = widthAdapter_1__T_63 | widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign widthAdapter_1__T_66 = ~widthAdapter_1__T_65; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign widthAdapter_1__T_67 = widthAdapter_1_ir0 == widthAdapter_1_ir4; // @[AXI4StreamWidthAdapter.scala 49:16]
  assign widthAdapter_1__T_69 = widthAdapter_1__T_67 | widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign widthAdapter_1__T_70 = ~widthAdapter_1__T_69; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign widthAdapter_1__GEN_6 = 2'h1 == widthAdapter_1__T_4 ? widthAdapter_1__T_1 : widthAdapter_1__T; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign widthAdapter_1_auto_in_ready = widthAdapter_1__T_6 & widthAdapter_1_auto_out_ready; // @[LazyModule.scala 173:31]
  assign widthAdapter_1_auto_out_valid = widthAdapter_1_auto_in_valid; // @[LazyModule.scala 173:49]
  assign widthAdapter_1_auto_out_bits_data = 2'h2 == widthAdapter_1__T_4 ? widthAdapter_1__T_2 : widthAdapter_1__GEN_6; // @[LazyModule.scala 173:49]
  assign widthAdapter_1_auto_out_bits_last = widthAdapter_1_auto_in_bits_last & widthAdapter_1__T_12; // @[LazyModule.scala 173:49]
  assign buffer_Queue__T_data__T_18_addr = buffer_Queue_value_1;
  assign buffer_Queue__T_data__T_18_data = buffer_Queue__T_data[buffer_Queue__T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_Queue__T_data__T_10_data = buffer_Queue_io_enq_bits_data;
  assign buffer_Queue__T_data__T_10_addr = buffer_Queue_value;
  assign buffer_Queue__T_data__T_10_mask = 1'h1;
  assign buffer_Queue__T_data__T_10_en = buffer_Queue_io_enq_ready & buffer_Queue_io_enq_valid;
  assign buffer_Queue__T_last__T_18_addr = buffer_Queue_value_1;
  assign buffer_Queue__T_last__T_18_data = buffer_Queue__T_last[buffer_Queue__T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_Queue__T_last__T_10_data = buffer_Queue_io_enq_bits_last;
  assign buffer_Queue__T_last__T_10_addr = buffer_Queue_value;
  assign buffer_Queue__T_last__T_10_mask = 1'h1;
  assign buffer_Queue__T_last__T_10_en = buffer_Queue_io_enq_ready & buffer_Queue_io_enq_valid;
  assign buffer_Queue__T_2 = buffer_Queue_value == buffer_Queue_value_1; // @[Decoupled.scala 214:41]
  assign buffer_Queue__T_3 = ~buffer_Queue__T_1; // @[Decoupled.scala 215:36]
  assign buffer_Queue__T_4 = buffer_Queue__T_2 & buffer_Queue__T_3; // @[Decoupled.scala 215:33]
  assign buffer_Queue__T_5 = buffer_Queue__T_2 & buffer_Queue__T_1; // @[Decoupled.scala 216:32]
  assign buffer_Queue__T_6 = buffer_Queue_io_enq_ready & buffer_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign buffer_Queue__T_8 = buffer_Queue_io_deq_ready & buffer_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign buffer_Queue__T_12 = buffer_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign buffer_Queue__T_14 = buffer_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign buffer_Queue__T_15 = buffer_Queue__T_6 != buffer_Queue__T_8; // @[Decoupled.scala 227:16]
  assign buffer_Queue_io_enq_ready = ~buffer_Queue__T_5; // @[Decoupled.scala 232:16]
  assign buffer_Queue_io_deq_valid = ~buffer_Queue__T_4; // @[Decoupled.scala 231:16]
  assign buffer_Queue_io_deq_bits_data = buffer_Queue__T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_Queue_io_deq_bits_last = buffer_Queue__T_last__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_auto_in_ready = buffer_Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign buffer_auto_out_valid = buffer_Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign buffer_auto_out_bits_data = buffer_Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign buffer_auto_out_bits_last = buffer_Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign buffer_Queue_clock = buffer_clock;
  assign buffer_Queue_reset = buffer_reset;
  assign buffer_Queue_io_enq_valid = buffer_auto_in_valid; // @[Decoupled.scala 288:22]
  assign buffer_Queue_io_enq_bits_data = buffer_auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign buffer_Queue_io_enq_bits_last = buffer_auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign buffer_Queue_io_deq_ready = buffer_auto_out_ready; // @[Decoupled.scala 311:15]
  assign buffer_1_Queue__T_data__T_18_addr = buffer_1_Queue_value_1;
  assign buffer_1_Queue__T_data__T_18_data = buffer_1_Queue__T_data[buffer_1_Queue__T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_1_Queue__T_data__T_10_data = buffer_1_Queue_io_enq_bits_data;
  assign buffer_1_Queue__T_data__T_10_addr = buffer_1_Queue_value;
  assign buffer_1_Queue__T_data__T_10_mask = 1'h1;
  assign buffer_1_Queue__T_data__T_10_en = buffer_1_Queue_io_enq_ready & buffer_1_Queue_io_enq_valid;
  assign buffer_1_Queue__T_last__T_18_addr = buffer_1_Queue_value_1;
  assign buffer_1_Queue__T_last__T_18_data = buffer_1_Queue__T_last[buffer_1_Queue__T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_1_Queue__T_last__T_10_data = buffer_1_Queue_io_enq_bits_last;
  assign buffer_1_Queue__T_last__T_10_addr = buffer_1_Queue_value;
  assign buffer_1_Queue__T_last__T_10_mask = 1'h1;
  assign buffer_1_Queue__T_last__T_10_en = buffer_1_Queue_io_enq_ready & buffer_1_Queue_io_enq_valid;
  assign buffer_1_Queue__T_2 = buffer_1_Queue_value == buffer_1_Queue_value_1; // @[Decoupled.scala 214:41]
  assign buffer_1_Queue__T_3 = ~buffer_1_Queue__T_1; // @[Decoupled.scala 215:36]
  assign buffer_1_Queue__T_4 = buffer_1_Queue__T_2 & buffer_1_Queue__T_3; // @[Decoupled.scala 215:33]
  assign buffer_1_Queue__T_5 = buffer_1_Queue__T_2 & buffer_1_Queue__T_1; // @[Decoupled.scala 216:32]
  assign buffer_1_Queue__T_6 = buffer_1_Queue_io_enq_ready & buffer_1_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign buffer_1_Queue__T_8 = buffer_1_Queue_io_deq_ready & buffer_1_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign buffer_1_Queue__T_12 = buffer_1_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign buffer_1_Queue__T_14 = buffer_1_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign buffer_1_Queue__T_15 = buffer_1_Queue__T_6 != buffer_1_Queue__T_8; // @[Decoupled.scala 227:16]
  assign buffer_1_Queue_io_enq_ready = ~buffer_1_Queue__T_5; // @[Decoupled.scala 232:16]
  assign buffer_1_Queue_io_deq_valid = ~buffer_1_Queue__T_4; // @[Decoupled.scala 231:16]
  assign buffer_1_Queue_io_deq_bits_data = buffer_1_Queue__T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_1_Queue_io_deq_bits_last = buffer_1_Queue__T_last__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_1_auto_in_ready = buffer_1_Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign buffer_1_auto_out_valid = buffer_1_Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign buffer_1_auto_out_bits_data = buffer_1_Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign buffer_1_auto_out_bits_last = buffer_1_Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign buffer_1_Queue_clock = buffer_1_clock;
  assign buffer_1_Queue_reset = buffer_1_reset;
  assign buffer_1_Queue_io_enq_valid = buffer_1_auto_in_valid; // @[Decoupled.scala 288:22]
  assign buffer_1_Queue_io_enq_bits_data = buffer_1_auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign buffer_1_Queue_io_enq_bits_last = buffer_1_auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign buffer_1_Queue_io_deq_ready = buffer_1_auto_out_ready; // @[Decoupled.scala 311:15]
  assign buffer_2_Queue__T_data__T_18_addr = buffer_2_Queue_value_1;
  assign buffer_2_Queue__T_data__T_18_data = buffer_2_Queue__T_data[buffer_2_Queue__T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_2_Queue__T_data__T_10_data = buffer_2_Queue_io_enq_bits_data;
  assign buffer_2_Queue__T_data__T_10_addr = buffer_2_Queue_value;
  assign buffer_2_Queue__T_data__T_10_mask = 1'h1;
  assign buffer_2_Queue__T_data__T_10_en = buffer_2_Queue_io_enq_ready & buffer_2_Queue_io_enq_valid;
  assign buffer_2_Queue__T_last__T_18_addr = buffer_2_Queue_value_1;
  assign buffer_2_Queue__T_last__T_18_data = buffer_2_Queue__T_last[buffer_2_Queue__T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_2_Queue__T_last__T_10_data = buffer_2_Queue_io_enq_bits_last;
  assign buffer_2_Queue__T_last__T_10_addr = buffer_2_Queue_value;
  assign buffer_2_Queue__T_last__T_10_mask = 1'h1;
  assign buffer_2_Queue__T_last__T_10_en = buffer_2_Queue_io_enq_ready & buffer_2_Queue_io_enq_valid;
  assign buffer_2_Queue__T_2 = buffer_2_Queue_value == buffer_2_Queue_value_1; // @[Decoupled.scala 214:41]
  assign buffer_2_Queue__T_3 = ~buffer_2_Queue__T_1; // @[Decoupled.scala 215:36]
  assign buffer_2_Queue__T_4 = buffer_2_Queue__T_2 & buffer_2_Queue__T_3; // @[Decoupled.scala 215:33]
  assign buffer_2_Queue__T_5 = buffer_2_Queue__T_2 & buffer_2_Queue__T_1; // @[Decoupled.scala 216:32]
  assign buffer_2_Queue__T_6 = buffer_2_Queue_io_enq_ready & buffer_2_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign buffer_2_Queue__T_8 = buffer_2_Queue_io_deq_ready & buffer_2_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign buffer_2_Queue__T_12 = buffer_2_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign buffer_2_Queue__T_14 = buffer_2_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign buffer_2_Queue__T_15 = buffer_2_Queue__T_6 != buffer_2_Queue__T_8; // @[Decoupled.scala 227:16]
  assign buffer_2_Queue_io_enq_ready = ~buffer_2_Queue__T_5; // @[Decoupled.scala 232:16]
  assign buffer_2_Queue_io_deq_valid = ~buffer_2_Queue__T_4; // @[Decoupled.scala 231:16]
  assign buffer_2_Queue_io_deq_bits_data = buffer_2_Queue__T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_2_Queue_io_deq_bits_last = buffer_2_Queue__T_last__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_2_auto_in_ready = buffer_2_Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign buffer_2_auto_out_valid = buffer_2_Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign buffer_2_auto_out_bits_data = buffer_2_Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign buffer_2_auto_out_bits_last = buffer_2_Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign buffer_2_Queue_clock = buffer_2_clock;
  assign buffer_2_Queue_reset = buffer_2_reset;
  assign buffer_2_Queue_io_enq_valid = buffer_2_auto_in_valid; // @[Decoupled.scala 288:22]
  assign buffer_2_Queue_io_enq_bits_data = buffer_2_auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign buffer_2_Queue_io_enq_bits_last = buffer_2_auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign buffer_2_Queue_io_deq_ready = buffer_2_auto_out_ready; // @[Decoupled.scala 311:15]
  assign buffer_3_Queue__T_data__T_18_addr = buffer_3_Queue_value_1;
  assign buffer_3_Queue__T_data__T_18_data = buffer_3_Queue__T_data[buffer_3_Queue__T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_3_Queue__T_data__T_10_data = buffer_3_Queue_io_enq_bits_data;
  assign buffer_3_Queue__T_data__T_10_addr = buffer_3_Queue_value;
  assign buffer_3_Queue__T_data__T_10_mask = 1'h1;
  assign buffer_3_Queue__T_data__T_10_en = buffer_3_Queue_io_enq_ready & buffer_3_Queue_io_enq_valid;
  assign buffer_3_Queue__T_last__T_18_addr = buffer_3_Queue_value_1;
  assign buffer_3_Queue__T_last__T_18_data = buffer_3_Queue__T_last[buffer_3_Queue__T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign buffer_3_Queue__T_last__T_10_data = buffer_3_Queue_io_enq_bits_last;
  assign buffer_3_Queue__T_last__T_10_addr = buffer_3_Queue_value;
  assign buffer_3_Queue__T_last__T_10_mask = 1'h1;
  assign buffer_3_Queue__T_last__T_10_en = buffer_3_Queue_io_enq_ready & buffer_3_Queue_io_enq_valid;
  assign buffer_3_Queue__T_2 = buffer_3_Queue_value == buffer_3_Queue_value_1; // @[Decoupled.scala 214:41]
  assign buffer_3_Queue__T_3 = ~buffer_3_Queue__T_1; // @[Decoupled.scala 215:36]
  assign buffer_3_Queue__T_4 = buffer_3_Queue__T_2 & buffer_3_Queue__T_3; // @[Decoupled.scala 215:33]
  assign buffer_3_Queue__T_5 = buffer_3_Queue__T_2 & buffer_3_Queue__T_1; // @[Decoupled.scala 216:32]
  assign buffer_3_Queue__T_6 = buffer_3_Queue_io_enq_ready & buffer_3_Queue_io_enq_valid; // @[Decoupled.scala 40:37]
  assign buffer_3_Queue__T_8 = buffer_3_Queue_io_deq_ready & buffer_3_Queue_io_deq_valid; // @[Decoupled.scala 40:37]
  assign buffer_3_Queue__T_12 = buffer_3_Queue_value + 1'h1; // @[Counter.scala 39:22]
  assign buffer_3_Queue__T_14 = buffer_3_Queue_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign buffer_3_Queue__T_15 = buffer_3_Queue__T_6 != buffer_3_Queue__T_8; // @[Decoupled.scala 227:16]
  assign buffer_3_Queue_io_enq_ready = ~buffer_3_Queue__T_5; // @[Decoupled.scala 232:16]
  assign buffer_3_Queue_io_deq_valid = ~buffer_3_Queue__T_4; // @[Decoupled.scala 231:16]
  assign buffer_3_Queue_io_deq_bits_data = buffer_3_Queue__T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_3_Queue_io_deq_bits_last = buffer_3_Queue__T_last__T_18_data; // @[Decoupled.scala 233:15]
  assign buffer_3_auto_in_ready = buffer_3_Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign buffer_3_auto_out_valid = buffer_3_Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign buffer_3_auto_out_bits_data = buffer_3_Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign buffer_3_auto_out_bits_last = buffer_3_Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign buffer_3_Queue_clock = buffer_3_clock;
  assign buffer_3_Queue_reset = buffer_3_reset;
  assign buffer_3_Queue_io_enq_valid = buffer_3_auto_in_valid; // @[Decoupled.scala 288:22]
  assign buffer_3_Queue_io_enq_bits_data = buffer_3_auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign buffer_3_Queue_io_enq_bits_last = buffer_3_auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign buffer_3_Queue_io_deq_ready = buffer_3_auto_out_ready; // @[Decoupled.scala 311:15]
  assign bus_awIn_0__T__T_18_addr = bus_awIn_0_value_1;
  assign bus_awIn_0__T__T_18_data = bus_awIn_0__T[bus_awIn_0__T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign bus_awIn_0__T__T_10_data = bus_awIn_0_io_enq_bits;
  assign bus_awIn_0__T__T_10_addr = bus_awIn_0_value;
  assign bus_awIn_0__T__T_10_mask = 1'h1;
  assign bus_awIn_0__T__T_10_en = bus_awIn_0__T_4 ? bus_awIn_0__GEN_9 : bus_awIn_0__T_6;
  assign bus_awIn_0__T_2 = bus_awIn_0_value == bus_awIn_0_value_1; // @[Decoupled.scala 214:41]
  assign bus_awIn_0__T_3 = ~bus_awIn_0__T_1; // @[Decoupled.scala 215:36]
  assign bus_awIn_0__T_4 = bus_awIn_0__T_2 & bus_awIn_0__T_3; // @[Decoupled.scala 215:33]
  assign bus_awIn_0__T_5 = bus_awIn_0__T_2 & bus_awIn_0__T_1; // @[Decoupled.scala 216:32]
  assign bus_awIn_0__T_6 = bus_awIn_0_io_enq_ready & bus_awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  assign bus_awIn_0__T_8 = bus_awIn_0_io_deq_ready & bus_awIn_0_io_deq_valid; // @[Decoupled.scala 40:37]
  assign bus_awIn_0__T_12 = bus_awIn_0_value + 1'h1; // @[Counter.scala 39:22]
  assign bus_awIn_0__GEN_9 = bus_awIn_0_io_deq_ready ? 1'h0 : bus_awIn_0__T_6; // @[Decoupled.scala 240:27]
  assign bus_awIn_0__GEN_12 = bus_awIn_0__T_4 ? bus_awIn_0__GEN_9 : bus_awIn_0__T_6; // @[Decoupled.scala 237:18]
  assign bus_awIn_0__T_14 = bus_awIn_0_value_1 + 1'h1; // @[Counter.scala 39:22]
  assign bus_awIn_0__GEN_11 = bus_awIn_0__T_4 ? 1'h0 : bus_awIn_0__T_8; // @[Decoupled.scala 237:18]
  assign bus_awIn_0__T_15 = bus_awIn_0__GEN_12 != bus_awIn_0__GEN_11; // @[Decoupled.scala 227:16]
  assign bus_awIn_0__T_16 = ~bus_awIn_0__T_4; // @[Decoupled.scala 231:19]
  assign bus_awIn_0_io_enq_ready = ~bus_awIn_0__T_5; // @[Decoupled.scala 232:16]
  assign bus_awIn_0_io_deq_valid = bus_awIn_0_io_enq_valid | bus_awIn_0__T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign bus_awIn_0_io_deq_bits = bus_awIn_0__T_4 ? bus_awIn_0_io_enq_bits : bus_awIn_0__T__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign bus__T_1 = {1'b0,$signed(bus_auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  assign bus__T_3 = $signed(bus__T_1) & 31'sh300; // @[Parameters.scala 137:52]
  assign bus_requestARIO_0_0 = $signed(bus__T_3) == 31'sh0; // @[Parameters.scala 137:67]
  assign bus__T_5 = bus_auto_in_ar_bits_addr ^ 30'h100; // @[Parameters.scala 137:31]
  assign bus__T_6 = {1'b0,$signed(bus__T_5)}; // @[Parameters.scala 137:49]
  assign bus__T_8 = $signed(bus__T_6) & 31'sh300; // @[Parameters.scala 137:52]
  assign bus_requestARIO_0_1 = $signed(bus__T_8) == 31'sh0; // @[Parameters.scala 137:67]
  assign bus__T_10 = bus_auto_in_ar_bits_addr ^ 30'h200; // @[Parameters.scala 137:31]
  assign bus__T_11 = {1'b0,$signed(bus__T_10)}; // @[Parameters.scala 137:49]
  assign bus__T_13 = $signed(bus__T_11) & 31'sh300; // @[Parameters.scala 137:52]
  assign bus_requestARIO_0_2 = $signed(bus__T_13) == 31'sh0; // @[Parameters.scala 137:67]
  assign bus__T_16 = {1'b0,$signed(bus_auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  assign bus__T_18 = $signed(bus__T_16) & 31'sh300; // @[Parameters.scala 137:52]
  assign bus_requestAWIO_0_0 = $signed(bus__T_18) == 31'sh0; // @[Parameters.scala 137:67]
  assign bus__T_20 = bus_auto_in_aw_bits_addr ^ 30'h100; // @[Parameters.scala 137:31]
  assign bus__T_21 = {1'b0,$signed(bus__T_20)}; // @[Parameters.scala 137:49]
  assign bus__T_23 = $signed(bus__T_21) & 31'sh300; // @[Parameters.scala 137:52]
  assign bus_requestAWIO_0_1 = $signed(bus__T_23) == 31'sh0; // @[Parameters.scala 137:67]
  assign bus__T_25 = bus_auto_in_aw_bits_addr ^ 30'h200; // @[Parameters.scala 137:31]
  assign bus__T_26 = {1'b0,$signed(bus__T_25)}; // @[Parameters.scala 137:49]
  assign bus__T_28 = $signed(bus__T_26) & 31'sh300; // @[Parameters.scala 137:52]
  assign bus_requestAWIO_0_2 = $signed(bus__T_28) == 31'sh0; // @[Parameters.scala 137:67]
  assign bus_requestROI_0_0 = ~bus_auto_out_0_r_bits_id; // @[Parameters.scala 47:9]
  assign bus_requestROI_1_0 = ~bus_auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  assign bus_requestROI_2_0 = ~bus_auto_out_2_r_bits_id; // @[Parameters.scala 47:9]
  assign bus_requestBOI_0_0 = ~bus_auto_out_0_b_bits_id; // @[Parameters.scala 47:9]
  assign bus_requestBOI_1_0 = ~bus_auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  assign bus_requestBOI_2_0 = ~bus_auto_out_2_b_bits_id; // @[Parameters.scala 47:9]
  assign bus__T_30 = {bus_requestAWIO_0_2,bus_requestAWIO_0_1}; // @[Xbar.scala 64:75]
  assign bus__T_31 = {bus_requestAWIO_0_2,bus_requestAWIO_0_1,bus_requestAWIO_0_0}; // @[Xbar.scala 64:75]
  assign bus_requestWIO_0_0 = bus_awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  assign bus_requestWIO_0_1 = bus_awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  assign bus_requestWIO_0_2 = bus_awIn_0_io_deq_bits[2]; // @[Xbar.scala 65:73]
  assign bus__T_39 = {bus_requestARIO_0_2,bus_requestARIO_0_1,bus_requestARIO_0_0}; // @[Xbar.scala 93:45]
  assign bus__T_40 = bus__T_39[2]; // @[OneHot.scala 30:18]
  assign bus__T_41 = bus__T_39[1:0]; // @[OneHot.scala 31:18]
  assign bus__GEN_22 = {{1'd0}, bus__T_40}; // @[OneHot.scala 32:28]
  assign bus__T_43 = bus__GEN_22 | bus__T_41; // @[OneHot.scala 32:28]
  assign bus__T_44 = bus__T_43[1]; // @[CircuitMath.scala 30:8]
  assign bus__T_45 = {bus__T_40,bus__T_44}; // @[Cat.scala 29:58]
  assign bus__T_48 = bus__T_31[2]; // @[OneHot.scala 30:18]
  assign bus__T_49 = bus__T_31[1:0]; // @[OneHot.scala 31:18]
  assign bus__GEN_23 = {{1'd0}, bus__T_48}; // @[OneHot.scala 32:28]
  assign bus__T_51 = bus__GEN_23 | bus__T_49; // @[OneHot.scala 32:28]
  assign bus__T_52 = bus__T_51[1]; // @[CircuitMath.scala 30:8]
  assign bus__T_53 = {bus__T_48,bus__T_52}; // @[Cat.scala 29:58]
  assign bus__T_132 = bus_requestARIO_0_0 & bus_auto_out_0_ar_ready; // @[Mux.scala 27:72]
  assign bus__T_133 = bus_requestARIO_0_1 & bus_auto_out_1_ar_ready; // @[Mux.scala 27:72]
  assign bus__T_135 = bus__T_132 | bus__T_133; // @[Mux.scala 27:72]
  assign bus__T_134 = bus_requestARIO_0_2 & bus_auto_out_2_ar_ready; // @[Mux.scala 27:72]
  assign bus_in_0_ar_ready = bus__T_135 | bus__T_134; // @[Mux.scala 27:72]
  assign bus__T_78 = bus__T_59 == 3'h0; // @[Xbar.scala 112:22]
  assign bus__T_77 = bus__T_60 == bus__T_45; // @[Xbar.scala 111:75]
  assign bus__T_79 = bus__T_78 | bus__T_77; // @[Xbar.scala 112:34]
  assign bus__T_80 = bus__T_59 != 3'h7; // @[Xbar.scala 112:80]
  assign bus__T_82 = bus__T_79 & bus__T_80; // @[Xbar.scala 112:48]
  assign bus_io_in_0_ar_ready = bus_in_0_ar_ready & bus__T_82; // @[Xbar.scala 130:45]
  assign bus__T_54 = bus_io_in_0_ar_ready & bus_auto_in_ar_valid; // @[Decoupled.scala 40:37]
  assign bus__T_159 = bus_auto_out_0_r_valid & bus_requestROI_0_0; // @[Xbar.scala 222:40]
  assign bus__T_161 = bus_auto_out_1_r_valid & bus_requestROI_1_0; // @[Xbar.scala 222:40]
  assign bus__T_303 = bus__T_159 | bus__T_161; // @[Xbar.scala 246:36]
  assign bus__T_163 = bus_auto_out_2_r_valid & bus_requestROI_2_0; // @[Xbar.scala 222:40]
  assign bus__T_304 = bus__T_303 | bus__T_163; // @[Xbar.scala 246:36]
  assign bus__T_380 = bus__T_373_0 & bus__T_159; // @[Mux.scala 27:72]
  assign bus__T_381 = bus__T_373_1 & bus__T_161; // @[Mux.scala 27:72]
  assign bus__T_383 = bus__T_380 | bus__T_381; // @[Mux.scala 27:72]
  assign bus__T_382 = bus__T_373_2 & bus__T_163; // @[Mux.scala 27:72]
  assign bus__T_384 = bus__T_383 | bus__T_382; // @[Mux.scala 27:72]
  assign bus_in_0_r_valid = bus__T_302 ? bus__T_304 : bus__T_384; // @[Xbar.scala 278:22]
  assign bus__T_56 = bus_auto_in_r_ready & bus_in_0_r_valid; // @[Decoupled.scala 40:37]
  assign bus__T_306 = {bus__T_163,bus__T_161,bus__T_159}; // @[Cat.scala 29:58]
  assign bus__T_314 = ~bus__T_313; // @[Arbiter.scala 21:30]
  assign bus__T_315 = bus__T_306 & bus__T_314; // @[Arbiter.scala 21:28]
  assign bus__T_316 = {bus__T_315,bus__T_163,bus__T_161,bus__T_159}; // @[Cat.scala 29:58]
  assign bus__T_317 = bus__T_316[5:1]; // @[package.scala 208:48]
  assign bus__GEN_24 = {{1'd0}, bus__T_317}; // @[package.scala 208:43]
  assign bus__T_318 = bus__T_316 | bus__GEN_24; // @[package.scala 208:43]
  assign bus__T_319 = bus__T_318[5:2]; // @[package.scala 208:48]
  assign bus__GEN_25 = {{2'd0}, bus__T_319}; // @[package.scala 208:43]
  assign bus__T_320 = bus__T_318 | bus__GEN_25; // @[package.scala 208:43]
  assign bus__T_322 = bus__T_320[5:1]; // @[Arbiter.scala 22:52]
  assign bus__T_323 = {bus__T_313, 3'h0}; // @[Arbiter.scala 22:66]
  assign bus__GEN_26 = {{1'd0}, bus__T_322}; // @[Arbiter.scala 22:58]
  assign bus__T_324 = bus__GEN_26 | bus__T_323; // @[Arbiter.scala 22:58]
  assign bus__T_325 = bus__T_324[5:3]; // @[Arbiter.scala 23:29]
  assign bus__T_326 = bus__T_324[2:0]; // @[Arbiter.scala 23:48]
  assign bus__T_327 = bus__T_325 & bus__T_326; // @[Arbiter.scala 23:39]
  assign bus__T_328 = ~bus__T_327; // @[Arbiter.scala 23:18]
  assign bus__T_340 = bus__T_328[0]; // @[Xbar.scala 248:69]
  assign bus__T_344 = bus__T_340 & bus__T_159; // @[Xbar.scala 250:63]
  assign bus__T_374_0 = bus__T_302 ? bus__T_344 : bus__T_373_0; // @[Xbar.scala 262:23]
  assign bus__T_389 = {bus_auto_out_0_r_bits_id,bus_auto_out_0_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  assign bus__T_390 = bus__T_374_0 ? bus__T_389 : 36'h0; // @[Mux.scala 27:72]
  assign bus__T_341 = bus__T_328[1]; // @[Xbar.scala 248:69]
  assign bus__T_345 = bus__T_341 & bus__T_161; // @[Xbar.scala 250:63]
  assign bus__T_374_1 = bus__T_302 ? bus__T_345 : bus__T_373_1; // @[Xbar.scala 262:23]
  assign bus__T_393 = {bus_auto_out_1_r_bits_id,bus_auto_out_1_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  assign bus__T_394 = bus__T_374_1 ? bus__T_393 : 36'h0; // @[Mux.scala 27:72]
  assign bus__T_399 = bus__T_390 | bus__T_394; // @[Mux.scala 27:72]
  assign bus__T_342 = bus__T_328[2]; // @[Xbar.scala 248:69]
  assign bus__T_346 = bus__T_342 & bus__T_163; // @[Xbar.scala 250:63]
  assign bus__T_374_2 = bus__T_302 ? bus__T_346 : bus__T_373_2; // @[Xbar.scala 262:23]
  assign bus__T_397 = {bus_auto_out_2_r_bits_id,bus_auto_out_2_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  assign bus__T_398 = bus__T_374_2 ? bus__T_397 : 36'h0; // @[Mux.scala 27:72]
  assign bus__T_400 = bus__T_399 | bus__T_398; // @[Mux.scala 27:72]
  assign bus_in_0_r_bits_last = bus__T_400[0]; // @[Mux.scala 27:72]
  assign bus__T_58 = bus__T_56 & bus_in_0_r_bits_last; // @[Xbar.scala 120:45]
  assign bus__GEN_27 = {{2'd0}, bus__T_54}; // @[Xbar.scala 106:30]
  assign bus__T_62 = bus__T_59 + bus__GEN_27; // @[Xbar.scala 106:30]
  assign bus__GEN_28 = {{2'd0}, bus__T_58}; // @[Xbar.scala 106:48]
  assign bus__T_64 = bus__T_62 - bus__GEN_28; // @[Xbar.scala 106:48]
  assign bus__T_65 = ~bus__T_58; // @[Xbar.scala 107:23]
  assign bus__T_66 = bus__T_59 != 3'h0; // @[Xbar.scala 107:43]
  assign bus__T_67 = bus__T_65 | bus__T_66; // @[Xbar.scala 107:34]
  assign bus__T_69 = bus__T_67 | bus_reset; // @[Xbar.scala 107:22]
  assign bus__T_70 = ~bus__T_69; // @[Xbar.scala 107:22]
  assign bus__T_71 = ~bus__T_54; // @[Xbar.scala 108:23]
  assign bus__T_73 = bus__T_71 | bus__T_80; // @[Xbar.scala 108:34]
  assign bus__T_75 = bus__T_73 | bus_reset; // @[Xbar.scala 108:22]
  assign bus__T_76 = ~bus__T_75; // @[Xbar.scala 108:22]
  assign bus__T_142 = bus_requestAWIO_0_0 & bus_auto_out_0_aw_ready; // @[Mux.scala 27:72]
  assign bus__T_143 = bus_requestAWIO_0_1 & bus_auto_out_1_aw_ready; // @[Mux.scala 27:72]
  assign bus__T_145 = bus__T_142 | bus__T_143; // @[Mux.scala 27:72]
  assign bus__T_144 = bus_requestAWIO_0_2 & bus_auto_out_2_aw_ready; // @[Mux.scala 27:72]
  assign bus_in_0_aw_ready = bus__T_145 | bus__T_144; // @[Mux.scala 27:72]
  assign bus__T_117 = bus__T_113 | bus_awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  assign bus__T_118 = bus_in_0_aw_ready & bus__T_117; // @[Xbar.scala 139:45]
  assign bus__T_106 = bus__T_87 == 3'h0; // @[Xbar.scala 112:22]
  assign bus__T_105 = bus__T_88 == bus__T_53; // @[Xbar.scala 111:75]
  assign bus__T_107 = bus__T_106 | bus__T_105; // @[Xbar.scala 112:34]
  assign bus__T_108 = bus__T_87 != 3'h7; // @[Xbar.scala 112:80]
  assign bus__T_110 = bus__T_107 & bus__T_108; // @[Xbar.scala 112:48]
  assign bus_io_in_0_aw_ready = bus__T_118 & bus__T_110; // @[Xbar.scala 139:82]
  assign bus__T_83 = bus_io_in_0_aw_ready & bus_auto_in_aw_valid; // @[Decoupled.scala 40:37]
  assign bus__T_165 = bus_auto_out_0_b_valid & bus_requestBOI_0_0; // @[Xbar.scala 222:40]
  assign bus__T_167 = bus_auto_out_1_b_valid & bus_requestBOI_1_0; // @[Xbar.scala 222:40]
  assign bus__T_408 = bus__T_165 | bus__T_167; // @[Xbar.scala 246:36]
  assign bus__T_169 = bus_auto_out_2_b_valid & bus_requestBOI_2_0; // @[Xbar.scala 222:40]
  assign bus__T_409 = bus__T_408 | bus__T_169; // @[Xbar.scala 246:36]
  assign bus__T_485 = bus__T_478_0 & bus__T_165; // @[Mux.scala 27:72]
  assign bus__T_486 = bus__T_478_1 & bus__T_167; // @[Mux.scala 27:72]
  assign bus__T_488 = bus__T_485 | bus__T_486; // @[Mux.scala 27:72]
  assign bus__T_487 = bus__T_478_2 & bus__T_169; // @[Mux.scala 27:72]
  assign bus__T_489 = bus__T_488 | bus__T_487; // @[Mux.scala 27:72]
  assign bus_in_0_b_valid = bus__T_407 ? bus__T_409 : bus__T_489; // @[Xbar.scala 278:22]
  assign bus__T_85 = bus_auto_in_b_ready & bus_in_0_b_valid; // @[Decoupled.scala 40:37]
  assign bus__GEN_29 = {{2'd0}, bus__T_83}; // @[Xbar.scala 106:30]
  assign bus__T_90 = bus__T_87 + bus__GEN_29; // @[Xbar.scala 106:30]
  assign bus__GEN_30 = {{2'd0}, bus__T_85}; // @[Xbar.scala 106:48]
  assign bus__T_92 = bus__T_90 - bus__GEN_30; // @[Xbar.scala 106:48]
  assign bus__T_93 = ~bus__T_85; // @[Xbar.scala 107:23]
  assign bus__T_94 = bus__T_87 != 3'h0; // @[Xbar.scala 107:43]
  assign bus__T_95 = bus__T_93 | bus__T_94; // @[Xbar.scala 107:34]
  assign bus__T_97 = bus__T_95 | bus_reset; // @[Xbar.scala 107:22]
  assign bus__T_98 = ~bus__T_97; // @[Xbar.scala 107:22]
  assign bus__T_99 = ~bus__T_83; // @[Xbar.scala 108:23]
  assign bus__T_101 = bus__T_99 | bus__T_108; // @[Xbar.scala 108:34]
  assign bus__T_103 = bus__T_101 | bus_reset; // @[Xbar.scala 108:22]
  assign bus__T_104 = ~bus__T_103; // @[Xbar.scala 108:22]
  assign bus_in_0_ar_valid = bus_auto_in_ar_valid & bus__T_82; // @[Xbar.scala 129:45]
  assign bus__T_115 = bus_auto_in_aw_valid & bus__T_117; // @[Xbar.scala 138:45]
  assign bus_in_0_aw_valid = bus__T_115 & bus__T_110; // @[Xbar.scala 138:82]
  assign bus__T_120 = ~bus__T_113; // @[Xbar.scala 140:54]
  assign bus__T_122 = bus_awIn_0_io_enq_ready & bus_awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  assign bus__GEN_2 = bus__T_122 | bus__T_113; // @[Xbar.scala 141:38]
  assign bus__T_123 = bus_in_0_aw_ready & bus_in_0_aw_valid; // @[Decoupled.scala 40:37]
  assign bus_in_0_w_valid = bus_auto_in_w_valid & bus_awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  assign bus__T_152 = bus_requestWIO_0_0 & bus_auto_out_0_w_ready; // @[Mux.scala 27:72]
  assign bus__T_153 = bus_requestWIO_0_1 & bus_auto_out_1_w_ready; // @[Mux.scala 27:72]
  assign bus__T_155 = bus__T_152 | bus__T_153; // @[Mux.scala 27:72]
  assign bus__T_154 = bus_requestWIO_0_2 & bus_auto_out_2_w_ready; // @[Mux.scala 27:72]
  assign bus_in_0_w_ready = bus__T_155 | bus__T_154; // @[Mux.scala 27:72]
  assign bus__T_126 = bus_auto_in_w_valid & bus_auto_in_w_bits_last; // @[Xbar.scala 147:50]
  assign bus_out_0_ar_valid = bus_in_0_ar_valid & bus_requestARIO_0_0; // @[Xbar.scala 222:40]
  assign bus_out_1_ar_valid = bus_in_0_ar_valid & bus_requestARIO_0_1; // @[Xbar.scala 222:40]
  assign bus_out_2_ar_valid = bus_in_0_ar_valid & bus_requestARIO_0_2; // @[Xbar.scala 222:40]
  assign bus_out_0_aw_valid = bus_in_0_aw_valid & bus_requestAWIO_0_0; // @[Xbar.scala 222:40]
  assign bus_out_1_aw_valid = bus_in_0_aw_valid & bus_requestAWIO_0_1; // @[Xbar.scala 222:40]
  assign bus_out_2_aw_valid = bus_in_0_aw_valid & bus_requestAWIO_0_2; // @[Xbar.scala 222:40]
  assign bus__T_176 = ~bus_out_0_aw_valid; // @[Xbar.scala 256:60]
  assign bus__T_182 = bus__T_176 | bus_out_0_aw_valid; // @[Xbar.scala 258:23]
  assign bus__T_184 = bus__T_182 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_185 = ~bus__T_184; // @[Xbar.scala 258:12]
  assign bus__T_197 = ~bus_out_0_ar_valid; // @[Xbar.scala 256:60]
  assign bus__T_203 = bus__T_197 | bus_out_0_ar_valid; // @[Xbar.scala 258:23]
  assign bus__T_205 = bus__T_203 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_206 = ~bus__T_205; // @[Xbar.scala 258:12]
  assign bus__T_220 = ~bus_out_1_aw_valid; // @[Xbar.scala 256:60]
  assign bus__T_226 = bus__T_220 | bus_out_1_aw_valid; // @[Xbar.scala 258:23]
  assign bus__T_228 = bus__T_226 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_229 = ~bus__T_228; // @[Xbar.scala 258:12]
  assign bus__T_241 = ~bus_out_1_ar_valid; // @[Xbar.scala 256:60]
  assign bus__T_247 = bus__T_241 | bus_out_1_ar_valid; // @[Xbar.scala 258:23]
  assign bus__T_249 = bus__T_247 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_250 = ~bus__T_249; // @[Xbar.scala 258:12]
  assign bus__T_264 = ~bus_out_2_aw_valid; // @[Xbar.scala 256:60]
  assign bus__T_270 = bus__T_264 | bus_out_2_aw_valid; // @[Xbar.scala 258:23]
  assign bus__T_272 = bus__T_270 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_273 = ~bus__T_272; // @[Xbar.scala 258:12]
  assign bus__T_285 = ~bus_out_2_ar_valid; // @[Xbar.scala 256:60]
  assign bus__T_291 = bus__T_285 | bus_out_2_ar_valid; // @[Xbar.scala 258:23]
  assign bus__T_293 = bus__T_291 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_294 = ~bus__T_293; // @[Xbar.scala 258:12]
  assign bus__T_329 = bus__T_306 != 3'h0; // @[Arbiter.scala 24:27]
  assign bus__T_330 = bus__T_302 & bus__T_329; // @[Arbiter.scala 24:18]
  assign bus__T_331 = bus__T_328 & bus__T_306; // @[Arbiter.scala 25:29]
  assign bus__T_332 = {bus__T_331, 1'h0}; // @[package.scala 199:48]
  assign bus__T_333 = bus__T_332[2:0]; // @[package.scala 199:53]
  assign bus__T_334 = bus__T_331 | bus__T_333; // @[package.scala 199:43]
  assign bus__T_335 = {bus__T_334, 2'h0}; // @[package.scala 199:48]
  assign bus__T_336 = bus__T_335[2:0]; // @[package.scala 199:53]
  assign bus__T_337 = bus__T_334 | bus__T_336; // @[package.scala 199:43]
  assign bus__T_349 = bus__T_344 | bus__T_345; // @[Xbar.scala 255:50]
  assign bus__T_350 = bus__T_349 | bus__T_346; // @[Xbar.scala 255:50]
  assign bus__T_352 = ~bus__T_344; // @[Xbar.scala 256:60]
  assign bus__T_355 = ~bus__T_345; // @[Xbar.scala 256:60]
  assign bus__T_356 = bus__T_352 | bus__T_355; // @[Xbar.scala 256:57]
  assign bus__T_357 = ~bus__T_349; // @[Xbar.scala 256:54]
  assign bus__T_358 = ~bus__T_346; // @[Xbar.scala 256:60]
  assign bus__T_359 = bus__T_357 | bus__T_358; // @[Xbar.scala 256:57]
  assign bus__T_361 = bus__T_356 & bus__T_359; // @[Xbar.scala 256:75]
  assign bus__T_363 = bus__T_361 | bus_reset; // @[Xbar.scala 256:11]
  assign bus__T_364 = ~bus__T_363; // @[Xbar.scala 256:11]
  assign bus__T_365 = ~bus__T_304; // @[Xbar.scala 258:13]
  assign bus__T_368 = bus__T_365 | bus__T_350; // @[Xbar.scala 258:23]
  assign bus__T_370 = bus__T_368 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_371 = ~bus__T_370; // @[Xbar.scala 258:12]
  assign bus__GEN_17 = bus__T_304 ? 1'h0 : bus__T_302; // @[Xbar.scala 266:21]
  assign bus__GEN_18 = bus__T_56 | bus__GEN_17; // @[Xbar.scala 267:24]
  assign bus__T_376_0 = bus__T_302 ? bus__T_340 : bus__T_373_0; // @[Xbar.scala 270:24]
  assign bus__T_376_1 = bus__T_302 ? bus__T_341 : bus__T_373_1; // @[Xbar.scala 270:24]
  assign bus__T_376_2 = bus__T_302 ? bus__T_342 : bus__T_373_2; // @[Xbar.scala 270:24]
  assign bus__T_411 = {bus__T_169,bus__T_167,bus__T_165}; // @[Cat.scala 29:58]
  assign bus__T_419 = ~bus__T_418; // @[Arbiter.scala 21:30]
  assign bus__T_420 = bus__T_411 & bus__T_419; // @[Arbiter.scala 21:28]
  assign bus__T_421 = {bus__T_420,bus__T_169,bus__T_167,bus__T_165}; // @[Cat.scala 29:58]
  assign bus__T_422 = bus__T_421[5:1]; // @[package.scala 208:48]
  assign bus__GEN_31 = {{1'd0}, bus__T_422}; // @[package.scala 208:43]
  assign bus__T_423 = bus__T_421 | bus__GEN_31; // @[package.scala 208:43]
  assign bus__T_424 = bus__T_423[5:2]; // @[package.scala 208:48]
  assign bus__GEN_32 = {{2'd0}, bus__T_424}; // @[package.scala 208:43]
  assign bus__T_425 = bus__T_423 | bus__GEN_32; // @[package.scala 208:43]
  assign bus__T_427 = bus__T_425[5:1]; // @[Arbiter.scala 22:52]
  assign bus__T_428 = {bus__T_418, 3'h0}; // @[Arbiter.scala 22:66]
  assign bus__GEN_33 = {{1'd0}, bus__T_427}; // @[Arbiter.scala 22:58]
  assign bus__T_429 = bus__GEN_33 | bus__T_428; // @[Arbiter.scala 22:58]
  assign bus__T_430 = bus__T_429[5:3]; // @[Arbiter.scala 23:29]
  assign bus__T_431 = bus__T_429[2:0]; // @[Arbiter.scala 23:48]
  assign bus__T_432 = bus__T_430 & bus__T_431; // @[Arbiter.scala 23:39]
  assign bus__T_433 = ~bus__T_432; // @[Arbiter.scala 23:18]
  assign bus__T_434 = bus__T_411 != 3'h0; // @[Arbiter.scala 24:27]
  assign bus__T_435 = bus__T_407 & bus__T_434; // @[Arbiter.scala 24:18]
  assign bus__T_436 = bus__T_433 & bus__T_411; // @[Arbiter.scala 25:29]
  assign bus__T_437 = {bus__T_436, 1'h0}; // @[package.scala 199:48]
  assign bus__T_438 = bus__T_437[2:0]; // @[package.scala 199:53]
  assign bus__T_439 = bus__T_436 | bus__T_438; // @[package.scala 199:43]
  assign bus__T_440 = {bus__T_439, 2'h0}; // @[package.scala 199:48]
  assign bus__T_441 = bus__T_440[2:0]; // @[package.scala 199:53]
  assign bus__T_442 = bus__T_439 | bus__T_441; // @[package.scala 199:43]
  assign bus__T_445 = bus__T_433[0]; // @[Xbar.scala 248:69]
  assign bus__T_446 = bus__T_433[1]; // @[Xbar.scala 248:69]
  assign bus__T_447 = bus__T_433[2]; // @[Xbar.scala 248:69]
  assign bus__T_449 = bus__T_445 & bus__T_165; // @[Xbar.scala 250:63]
  assign bus__T_450 = bus__T_446 & bus__T_167; // @[Xbar.scala 250:63]
  assign bus__T_451 = bus__T_447 & bus__T_169; // @[Xbar.scala 250:63]
  assign bus__T_454 = bus__T_449 | bus__T_450; // @[Xbar.scala 255:50]
  assign bus__T_455 = bus__T_454 | bus__T_451; // @[Xbar.scala 255:50]
  assign bus__T_457 = ~bus__T_449; // @[Xbar.scala 256:60]
  assign bus__T_460 = ~bus__T_450; // @[Xbar.scala 256:60]
  assign bus__T_461 = bus__T_457 | bus__T_460; // @[Xbar.scala 256:57]
  assign bus__T_462 = ~bus__T_454; // @[Xbar.scala 256:54]
  assign bus__T_463 = ~bus__T_451; // @[Xbar.scala 256:60]
  assign bus__T_464 = bus__T_462 | bus__T_463; // @[Xbar.scala 256:57]
  assign bus__T_466 = bus__T_461 & bus__T_464; // @[Xbar.scala 256:75]
  assign bus__T_468 = bus__T_466 | bus_reset; // @[Xbar.scala 256:11]
  assign bus__T_469 = ~bus__T_468; // @[Xbar.scala 256:11]
  assign bus__T_470 = ~bus__T_409; // @[Xbar.scala 258:13]
  assign bus__T_473 = bus__T_470 | bus__T_455; // @[Xbar.scala 258:23]
  assign bus__T_475 = bus__T_473 | bus_reset; // @[Xbar.scala 258:12]
  assign bus__T_476 = ~bus__T_475; // @[Xbar.scala 258:12]
  assign bus__T_479_0 = bus__T_407 ? bus__T_449 : bus__T_478_0; // @[Xbar.scala 262:23]
  assign bus__T_479_1 = bus__T_407 ? bus__T_450 : bus__T_478_1; // @[Xbar.scala 262:23]
  assign bus__T_479_2 = bus__T_407 ? bus__T_451 : bus__T_478_2; // @[Xbar.scala 262:23]
  assign bus__GEN_20 = bus__T_409 ? 1'h0 : bus__T_407; // @[Xbar.scala 266:21]
  assign bus__GEN_21 = bus__T_85 | bus__GEN_20; // @[Xbar.scala 267:24]
  assign bus__T_481_0 = bus__T_407 ? bus__T_445 : bus__T_478_0; // @[Xbar.scala 270:24]
  assign bus__T_481_1 = bus__T_407 ? bus__T_446 : bus__T_478_1; // @[Xbar.scala 270:24]
  assign bus__T_481_2 = bus__T_407 ? bus__T_447 : bus__T_478_2; // @[Xbar.scala 270:24]
  assign bus__T_492 = {bus_auto_out_0_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  assign bus__T_493 = bus__T_479_0 ? bus__T_492 : 3'h0; // @[Mux.scala 27:72]
  assign bus__T_494 = {bus_auto_out_1_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  assign bus__T_495 = bus__T_479_1 ? bus__T_494 : 3'h0; // @[Mux.scala 27:72]
  assign bus__T_496 = {bus_auto_out_2_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  assign bus__T_497 = bus__T_479_2 ? bus__T_496 : 3'h0; // @[Mux.scala 27:72]
  assign bus__T_498 = bus__T_493 | bus__T_495; // @[Mux.scala 27:72]
  assign bus__T_499 = bus__T_498 | bus__T_497; // @[Mux.scala 27:72]
  assign bus_auto_in_aw_ready = bus__T_118 & bus__T_110; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_ready = bus_in_0_w_ready & bus_awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign bus_auto_in_b_valid = bus__T_407 ? bus__T_409 : bus__T_489; // @[LazyModule.scala 173:31]
  assign bus_auto_in_b_bits_resp = bus__T_499[1:0]; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_ready = bus_in_0_ar_ready & bus__T_82; // @[LazyModule.scala 173:31]
  assign bus_auto_in_r_valid = bus__T_302 ? bus__T_304 : bus__T_384; // @[LazyModule.scala 173:31]
  assign bus_auto_in_r_bits_data = bus__T_400[34:3]; // @[LazyModule.scala 173:31]
  assign bus_auto_in_r_bits_resp = bus__T_400[2:1]; // @[LazyModule.scala 173:31]
  assign bus_auto_in_r_bits_last = bus__T_400[0]; // @[LazyModule.scala 173:31]
  assign bus_auto_out_2_aw_valid = bus_in_0_aw_valid & bus_requestAWIO_0_2; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_aw_bits_id = bus_auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_aw_bits_addr = bus_auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_w_valid = bus_in_0_w_valid & bus_requestWIO_0_2; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_w_bits_data = bus_auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_w_bits_strb = bus_auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_b_ready = bus_auto_in_b_ready & bus__T_481_2; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_ar_valid = bus_in_0_ar_valid & bus_requestARIO_0_2; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_ar_bits_id = bus_auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_ar_bits_addr = bus_auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_ar_bits_size = bus_auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign bus_auto_out_2_r_ready = bus_auto_in_r_ready & bus__T_376_2; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_aw_valid = bus_in_0_aw_valid & bus_requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_aw_bits_id = bus_auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_aw_bits_addr = bus_auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_w_valid = bus_in_0_w_valid & bus_requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_w_bits_data = bus_auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_w_bits_strb = bus_auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_b_ready = bus_auto_in_b_ready & bus__T_481_1; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_ar_valid = bus_in_0_ar_valid & bus_requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_ar_bits_id = bus_auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_ar_bits_addr = bus_auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_ar_bits_size = bus_auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign bus_auto_out_1_r_ready = bus_auto_in_r_ready & bus__T_376_1; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_aw_valid = bus_in_0_aw_valid & bus_requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_aw_bits_id = bus_auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_aw_bits_addr = bus_auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_w_valid = bus_in_0_w_valid & bus_requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_b_ready = bus_auto_in_b_ready & bus__T_481_0; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_ar_valid = bus_in_0_ar_valid & bus_requestARIO_0_0; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_ar_bits_id = bus_auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_ar_bits_addr = bus_auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign bus_auto_out_0_r_ready = bus_auto_in_r_ready & bus__T_376_0; // @[LazyModule.scala 173:49]
  assign bus_awIn_0_clock = bus_clock;
  assign bus_awIn_0_reset = bus_reset;
  assign bus_awIn_0_io_enq_valid = bus_auto_in_aw_valid & bus__T_120; // @[Xbar.scala 140:30]
  assign bus_awIn_0_io_enq_bits = {bus__T_30,bus_requestAWIO_0_0}; // @[Xbar.scala 64:57]
  assign bus_awIn_0_io_deq_ready = bus__T_126 & bus_in_0_w_ready; // @[Xbar.scala 147:30]
  assign converter_auto_in_aw_ready = converter_auto_out_aw_ready; // @[LazyModule.scala 173:31]
  assign converter_auto_in_w_ready = converter_auto_out_w_ready; // @[LazyModule.scala 173:31]
  assign converter_auto_in_b_valid = converter_auto_out_b_valid; // @[LazyModule.scala 173:31]
  assign converter_auto_in_b_bits_resp = converter_auto_out_b_bits_resp; // @[LazyModule.scala 173:31]
  assign converter_auto_in_ar_ready = converter_auto_out_ar_ready; // @[LazyModule.scala 173:31]
  assign converter_auto_in_r_valid = converter_auto_out_r_valid; // @[LazyModule.scala 173:31]
  assign converter_auto_in_r_bits_data = converter_auto_out_r_bits_data; // @[LazyModule.scala 173:31]
  assign converter_auto_in_r_bits_resp = converter_auto_out_r_bits_resp; // @[LazyModule.scala 173:31]
  assign converter_auto_in_r_bits_last = converter_auto_out_r_bits_last; // @[LazyModule.scala 173:31]
  assign converter_auto_out_aw_valid = converter_auto_in_aw_valid; // @[LazyModule.scala 173:49]
  assign converter_auto_out_aw_bits_id = converter_auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign converter_auto_out_aw_bits_addr = converter_auto_in_aw_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign converter_auto_out_w_valid = converter_auto_in_w_valid; // @[LazyModule.scala 173:49]
  assign converter_auto_out_w_bits_data = converter_auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign converter_auto_out_w_bits_strb = converter_auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign converter_auto_out_w_bits_last = converter_auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign converter_auto_out_b_ready = converter_auto_in_b_ready; // @[LazyModule.scala 173:49]
  assign converter_auto_out_ar_valid = converter_auto_in_ar_valid; // @[LazyModule.scala 173:49]
  assign converter_auto_out_ar_bits_id = converter_auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign converter_auto_out_ar_bits_addr = converter_auto_in_ar_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign converter_auto_out_ar_bits_size = converter_auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign converter_auto_out_r_ready = converter_auto_in_r_ready; // @[LazyModule.scala 173:49]
  assign converter_1_auto_in_ready = converter_1_auto_out_ready; // @[LazyModule.scala 173:31]
  assign converter_1_auto_out_valid = converter_1_auto_in_valid; // @[LazyModule.scala 173:49]
  assign converter_1_auto_out_bits_data = converter_1_auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign converter_1_auto_out_bits_last = converter_1_auto_in_bits_last; // @[LazyModule.scala 173:49]
  assign converter_2_auto_in_ready = converter_2_auto_out_ready; // @[LazyModule.scala 173:31]
  assign converter_2_auto_out_valid = converter_2_auto_in_valid; // @[LazyModule.scala 173:49]
  assign converter_2_auto_out_bits_data = converter_2_auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign converter_2_auto_out_bits_last = converter_2_auto_in_bits_last; // @[LazyModule.scala 173:49]
  assign ioMem_0_aw_ready = converter_auto_in_aw_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_w_ready = converter_auto_in_w_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_b_valid = converter_auto_in_b_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_resp = converter_auto_in_b_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_ar_ready = converter_auto_in_ar_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_r_valid = converter_auto_in_r_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_data = converter_auto_in_r_bits_data; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_resp = converter_auto_in_r_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_last = converter_auto_in_r_bits_last; // @[Nodes.scala 624:60]
  assign in_0_ready = converter_2_auto_in_ready; // @[Nodes.scala 624:60]
  assign out_0_valid = converter_1_auto_out_valid; // @[Nodes.scala 649:56]
  assign out_0_bits_data = converter_1_auto_out_bits_data; // @[Nodes.scala 649:56]
  assign out_0_bits_last = converter_1_auto_out_bits_last; // @[Nodes.scala 649:56]
  assign widthAdapter_clock = clock;
  assign widthAdapter_reset = reset;
  assign widthAdapter_auto_in_valid = converter_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_data = converter_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_last = converter_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_out_ready = buffer_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_auto_mem_in_aw_valid = bus_auto_out_0_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_id = bus_auto_out_0_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_addr = bus_auto_out_0_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_valid = bus_auto_out_0_w_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_b_ready = bus_auto_out_0_b_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_valid = bus_auto_out_0_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_id = bus_auto_out_0_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_addr = bus_auto_out_0_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_r_ready = bus_auto_out_0_r_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_valid = buffer_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_data = buffer_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_last = buffer_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_out_ready = buffer_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_clock = clock;
  assign mag_reset = reset;
  assign mag_auto_mem_in_aw_valid = bus_auto_out_1_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_id = bus_auto_out_1_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_addr = bus_auto_out_1_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_valid = bus_auto_out_1_w_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_data = bus_auto_out_1_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_strb = bus_auto_out_1_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_b_ready = bus_auto_out_1_b_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_valid = bus_auto_out_1_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_id = bus_auto_out_1_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_addr = bus_auto_out_1_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_size = bus_auto_out_1_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_r_ready = bus_auto_out_1_r_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_master_out_ready = buffer_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_auto_slave_in_valid = buffer_auto_out_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_slave_in_bits_data = buffer_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_slave_in_bits_last = buffer_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign cfar_clock = clock;
  assign cfar_reset = reset;
  assign cfar_auto_mem_in_aw_valid = bus_auto_out_2_aw_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_aw_bits_id = bus_auto_out_2_aw_bits_id; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_aw_bits_addr = bus_auto_out_2_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_w_valid = bus_auto_out_2_w_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_w_bits_data = bus_auto_out_2_w_bits_data; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_w_bits_strb = bus_auto_out_2_w_bits_strb; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_b_ready = bus_auto_out_2_b_ready; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_valid = bus_auto_out_2_ar_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_bits_id = bus_auto_out_2_ar_bits_id; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_bits_addr = bus_auto_out_2_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_bits_size = bus_auto_out_2_ar_bits_size; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_r_ready = bus_auto_out_2_r_ready; // @[LazyModule.scala 167:31]
  assign cfar_auto_master_out_ready = buffer_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign cfar_auto_slave_in_valid = buffer_1_auto_out_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_slave_in_bits_data = buffer_1_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign cfar_auto_slave_in_bits_last = buffer_1_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_clock = clock;
  assign widthAdapter_1_reset = reset;
  assign widthAdapter_1_auto_in_valid = buffer_3_auto_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_auto_in_bits_data = buffer_3_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_auto_in_bits_last = buffer_3_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_auto_out_ready = converter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_valid = fft_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_data = fft_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_last = fft_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_auto_out_ready = mag_auto_slave_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_1_clock = clock;
  assign buffer_1_reset = reset;
  assign buffer_1_auto_in_valid = mag_auto_master_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_data = mag_auto_master_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_last = mag_auto_master_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_out_ready = cfar_auto_slave_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_2_clock = clock;
  assign buffer_2_reset = reset;
  assign buffer_2_auto_in_valid = widthAdapter_auto_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_data = widthAdapter_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_last = widthAdapter_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_out_ready = fft_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_3_clock = clock;
  assign buffer_3_reset = reset;
  assign buffer_3_auto_in_valid = cfar_auto_master_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_data = cfar_auto_master_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_last = cfar_auto_master_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_out_ready = widthAdapter_1_auto_in_ready; // @[LazyModule.scala 167:31]
  assign bus_clock = clock;
  assign bus_reset = reset;
  assign bus_auto_in_aw_valid = converter_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_id = converter_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_addr = converter_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_valid = converter_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_data = converter_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_strb = converter_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_last = converter_auto_out_w_bits_last; // @[LazyModule.scala 167:31]
  assign bus_auto_in_b_ready = converter_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_valid = converter_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_id = converter_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_addr = converter_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_size = converter_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_r_ready = converter_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_aw_ready = cfar_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_w_ready = cfar_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_b_valid = cfar_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_b_bits_id = cfar_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_ar_ready = cfar_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_r_valid = cfar_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_r_bits_id = cfar_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_r_bits_data = cfar_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_aw_ready = mag_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_w_ready = mag_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_b_valid = mag_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_b_bits_id = mag_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_ar_ready = mag_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_r_valid = mag_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_r_bits_id = mag_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_r_bits_data = mag_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_aw_ready = fft_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_w_ready = fft_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_b_valid = fft_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_b_bits_id = fft_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_ar_ready = fft_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_r_valid = fft_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_r_bits_id = fft_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_r_bits_data = fft_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign converter_auto_in_aw_valid = ioMem_0_aw_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_id = ioMem_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_addr = ioMem_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_valid = ioMem_0_w_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_data = ioMem_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_strb = ioMem_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_last = ioMem_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign converter_auto_in_b_ready = ioMem_0_b_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_valid = ioMem_0_ar_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_id = ioMem_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_addr = ioMem_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_size = ioMem_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_r_ready = ioMem_0_r_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_out_aw_ready = bus_auto_in_aw_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_w_ready = bus_auto_in_w_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_valid = bus_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_bits_resp = bus_auto_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_ar_ready = bus_auto_in_ar_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_valid = bus_auto_in_r_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_data = bus_auto_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_resp = bus_auto_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_last = bus_auto_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign converter_1_auto_in_valid = widthAdapter_1_auto_out_valid; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_data = widthAdapter_1_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_last = widthAdapter_1_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign converter_1_auto_out_ready = out_0_ready; // @[LazyModule.scala 167:31]
  assign converter_2_auto_in_valid = in_0_valid; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_data = in_0_bits_data; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_last = in_0_bits_last; // @[LazyModule.scala 167:57]
  assign converter_2_auto_out_ready = widthAdapter_auto_in_ready; // @[LazyModule.scala 167:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  widthAdapter__T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  widthAdapter__T_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  widthAdapter__T_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  widthAdapter__T_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  widthAdapter__T_20 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  widthAdapter__T_21 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  widthAdapter__T_22 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  widthAdapter__T_23 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  widthAdapter__T_44 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  widthAdapter__T_64 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  widthAdapter__T_84 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_0_feedback_real = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_0_feedback_imag = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_1_feedback_real = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_1_feedback_imag = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_1__T_21_real = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_1__T_21_imag = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2_feedback_real = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2_feedback_imag = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2__T_21_real = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2__T_21_imag = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2__T_24_real = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2__T_24_imag = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2__T_27_real = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_2__T_27_imag = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3_feedback_real = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3_feedback_imag = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_21_real = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_21_imag = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_24_real = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_24_imag = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_27_real = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_27_imag = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_30_real = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_30_imag = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_33_real = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_33_imag = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_36_real = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_36_imag = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_39_real = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_3__T_39_imag = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4_feedback_real = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4_feedback_imag = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_21_real = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_21_imag = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_24_real = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_24_imag = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_27_real = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_27_imag = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_30_real = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_30_imag = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_33_real = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_33_imag = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_36_real = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_36_imag = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_39_real = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_39_imag = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_42_real = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_42_imag = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_45_real = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_45_imag = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_48_real = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_48_imag = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_51_real = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_51_imag = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_54_real = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_54_imag = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_57_real = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_57_imag = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_60_real = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_60_imag = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_63_real = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_4__T_63_imag = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5_feedback_real = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5_feedback_imag = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_21_real = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_21_imag = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_24_real = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_24_imag = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_27_real = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_27_imag = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_30_real = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_30_imag = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_33_real = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_33_imag = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_36_real = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_36_imag = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_39_real = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_39_imag = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_42_real = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_42_imag = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_45_real = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_45_imag = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_48_real = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_48_imag = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_51_real = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_51_imag = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_54_real = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_54_imag = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_57_real = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_57_imag = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_60_real = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_60_imag = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_63_real = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_63_imag = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_66_real = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_66_imag = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_69_real = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_69_imag = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_72_real = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_72_imag = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_75_real = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_75_imag = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_78_real = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_78_imag = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_81_real = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_81_imag = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_84_real = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_84_imag = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_87_real = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_87_imag = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_90_real = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_90_imag = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_93_real = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_93_imag = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_96_real = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_96_imag = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_99_real = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_99_imag = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_102_real = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_102_imag = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_105_real = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_105_imag = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_108_real = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_108_imag = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_111_real = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_5__T_111_imag = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6_feedback_real = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6_feedback_imag = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_21_real = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_21_imag = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_24_real = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_24_imag = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_27_real = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_27_imag = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_30_real = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_30_imag = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_33_real = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_33_imag = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_36_real = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_36_imag = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_39_real = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_39_imag = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_42_real = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_42_imag = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_45_real = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_45_imag = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_48_real = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_48_imag = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_51_real = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_51_imag = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_54_real = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_54_imag = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_57_real = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_57_imag = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_60_real = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_60_imag = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_63_real = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_63_imag = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_66_real = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_66_imag = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_69_real = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_69_imag = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_72_real = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_72_imag = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_75_real = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_75_imag = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_78_real = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_78_imag = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_81_real = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_81_imag = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_84_real = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_84_imag = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_87_real = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_87_imag = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_90_real = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_90_imag = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_93_real = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_93_imag = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_96_real = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_96_imag = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_99_real = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_99_imag = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_102_real = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_102_imag = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_105_real = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_105_imag = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_108_real = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_108_imag = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_111_real = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_111_imag = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_114_real = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_114_imag = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_117_real = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_117_imag = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_120_real = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_120_imag = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_123_real = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_123_imag = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_126_real = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_126_imag = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_129_real = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_129_imag = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_132_real = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_132_imag = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_135_real = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_135_imag = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_138_real = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_138_imag = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_141_real = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_141_imag = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_144_real = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_144_imag = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_147_real = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_147_imag = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_150_real = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_150_imag = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_153_real = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_153_imag = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_156_real = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_156_imag = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_159_real = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_159_imag = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_162_real = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_162_imag = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_165_real = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_165_imag = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_168_real = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_168_imag = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_171_real = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_171_imag = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_174_real = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_174_imag = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_177_real = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_177_imag = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_180_real = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_180_imag = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_183_real = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_183_imag = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_186_real = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_186_imag = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_189_real = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_189_imag = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_192_real = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_192_imag = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_195_real = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_195_imag = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_198_real = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_198_imag = _RAND_258[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_201_real = _RAND_259[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_201_imag = _RAND_260[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_204_real = _RAND_261[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_204_imag = _RAND_262[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_207_real = _RAND_263[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_6__T_207_imag = _RAND_264[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7_feedback_real = _RAND_265[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7_feedback_imag = _RAND_266[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_21_real = _RAND_267[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_21_imag = _RAND_268[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_24_real = _RAND_269[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_24_imag = _RAND_270[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_27_real = _RAND_271[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_27_imag = _RAND_272[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_30_real = _RAND_273[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_30_imag = _RAND_274[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_33_real = _RAND_275[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_33_imag = _RAND_276[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_36_real = _RAND_277[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_36_imag = _RAND_278[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_39_real = _RAND_279[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_39_imag = _RAND_280[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_42_real = _RAND_281[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_42_imag = _RAND_282[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_45_real = _RAND_283[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_45_imag = _RAND_284[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_48_real = _RAND_285[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_48_imag = _RAND_286[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_51_real = _RAND_287[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_51_imag = _RAND_288[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_54_real = _RAND_289[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_54_imag = _RAND_290[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_57_real = _RAND_291[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_57_imag = _RAND_292[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_60_real = _RAND_293[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_60_imag = _RAND_294[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_63_real = _RAND_295[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_63_imag = _RAND_296[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_66_real = _RAND_297[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_66_imag = _RAND_298[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_69_real = _RAND_299[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_69_imag = _RAND_300[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_72_real = _RAND_301[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_72_imag = _RAND_302[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_75_real = _RAND_303[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_75_imag = _RAND_304[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_78_real = _RAND_305[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_78_imag = _RAND_306[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_81_real = _RAND_307[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_81_imag = _RAND_308[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_84_real = _RAND_309[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_84_imag = _RAND_310[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_87_real = _RAND_311[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_87_imag = _RAND_312[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_90_real = _RAND_313[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_90_imag = _RAND_314[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_93_real = _RAND_315[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_93_imag = _RAND_316[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_96_real = _RAND_317[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_96_imag = _RAND_318[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_99_real = _RAND_319[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_99_imag = _RAND_320[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_102_real = _RAND_321[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_102_imag = _RAND_322[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_105_real = _RAND_323[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_105_imag = _RAND_324[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_108_real = _RAND_325[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_108_imag = _RAND_326[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_111_real = _RAND_327[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_111_imag = _RAND_328[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_114_real = _RAND_329[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_114_imag = _RAND_330[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_117_real = _RAND_331[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_117_imag = _RAND_332[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_120_real = _RAND_333[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_120_imag = _RAND_334[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_123_real = _RAND_335[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_123_imag = _RAND_336[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_126_real = _RAND_337[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_126_imag = _RAND_338[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_129_real = _RAND_339[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_129_imag = _RAND_340[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_132_real = _RAND_341[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_132_imag = _RAND_342[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_135_real = _RAND_343[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_135_imag = _RAND_344[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_138_real = _RAND_345[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_138_imag = _RAND_346[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_141_real = _RAND_347[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_141_imag = _RAND_348[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_144_real = _RAND_349[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_144_imag = _RAND_350[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_147_real = _RAND_351[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_147_imag = _RAND_352[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_150_real = _RAND_353[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_150_imag = _RAND_354[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_153_real = _RAND_355[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_153_imag = _RAND_356[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_156_real = _RAND_357[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_156_imag = _RAND_358[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_159_real = _RAND_359[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_159_imag = _RAND_360[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_162_real = _RAND_361[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_162_imag = _RAND_362[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_165_real = _RAND_363[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_165_imag = _RAND_364[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_168_real = _RAND_365[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_168_imag = _RAND_366[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_171_real = _RAND_367[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_171_imag = _RAND_368[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_174_real = _RAND_369[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_174_imag = _RAND_370[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_177_real = _RAND_371[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_177_imag = _RAND_372[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_180_real = _RAND_373[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_180_imag = _RAND_374[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_183_real = _RAND_375[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_183_imag = _RAND_376[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_186_real = _RAND_377[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_186_imag = _RAND_378[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_189_real = _RAND_379[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_189_imag = _RAND_380[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_192_real = _RAND_381[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_192_imag = _RAND_382[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_195_real = _RAND_383[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_195_imag = _RAND_384[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_198_real = _RAND_385[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_198_imag = _RAND_386[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_201_real = _RAND_387[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_201_imag = _RAND_388[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_204_real = _RAND_389[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_204_imag = _RAND_390[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_207_real = _RAND_391[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_207_imag = _RAND_392[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_210_real = _RAND_393[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_210_imag = _RAND_394[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_213_real = _RAND_395[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_213_imag = _RAND_396[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_216_real = _RAND_397[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_216_imag = _RAND_398[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_219_real = _RAND_399[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_219_imag = _RAND_400[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_222_real = _RAND_401[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_222_imag = _RAND_402[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_225_real = _RAND_403[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_225_imag = _RAND_404[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_228_real = _RAND_405[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_228_imag = _RAND_406[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_231_real = _RAND_407[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_231_imag = _RAND_408[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_234_real = _RAND_409[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_234_imag = _RAND_410[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_237_real = _RAND_411[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_237_imag = _RAND_412[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_240_real = _RAND_413[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_240_imag = _RAND_414[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_243_real = _RAND_415[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_243_imag = _RAND_416[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_246_real = _RAND_417[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_246_imag = _RAND_418[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_249_real = _RAND_419[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_249_imag = _RAND_420[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_252_real = _RAND_421[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_252_imag = _RAND_422[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_255_real = _RAND_423[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_255_imag = _RAND_424[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_258_real = _RAND_425[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_258_imag = _RAND_426[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_261_real = _RAND_427[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_261_imag = _RAND_428[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_264_real = _RAND_429[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_264_imag = _RAND_430[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_267_real = _RAND_431[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_267_imag = _RAND_432[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_270_real = _RAND_433[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_270_imag = _RAND_434[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_273_real = _RAND_435[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_273_imag = _RAND_436[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_276_real = _RAND_437[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_276_imag = _RAND_438[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_279_real = _RAND_439[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_279_imag = _RAND_440[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_282_real = _RAND_441[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_282_imag = _RAND_442[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_285_real = _RAND_443[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_285_imag = _RAND_444[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_288_real = _RAND_445[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_288_imag = _RAND_446[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_291_real = _RAND_447[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_291_imag = _RAND_448[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_294_real = _RAND_449[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_294_imag = _RAND_450[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_297_real = _RAND_451[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_297_imag = _RAND_452[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_300_real = _RAND_453[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_300_imag = _RAND_454[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_303_real = _RAND_455[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_303_imag = _RAND_456[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_306_real = _RAND_457[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_306_imag = _RAND_458[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_309_real = _RAND_459[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_309_imag = _RAND_460[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_312_real = _RAND_461[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_312_imag = _RAND_462[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_315_real = _RAND_463[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_315_imag = _RAND_464[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_318_real = _RAND_465[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_318_imag = _RAND_466[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_321_real = _RAND_467[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_321_imag = _RAND_468[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_324_real = _RAND_469[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_324_imag = _RAND_470[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_327_real = _RAND_471[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_327_imag = _RAND_472[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_330_real = _RAND_473[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_330_imag = _RAND_474[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_333_real = _RAND_475[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_333_imag = _RAND_476[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_336_real = _RAND_477[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_336_imag = _RAND_478[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_339_real = _RAND_479[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_339_imag = _RAND_480[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_342_real = _RAND_481[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_342_imag = _RAND_482[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_345_real = _RAND_483[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_345_imag = _RAND_484[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_348_real = _RAND_485[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_348_imag = _RAND_486[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_351_real = _RAND_487[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_351_imag = _RAND_488[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_354_real = _RAND_489[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_354_imag = _RAND_490[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_357_real = _RAND_491[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_357_imag = _RAND_492[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_360_real = _RAND_493[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_360_imag = _RAND_494[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_363_real = _RAND_495[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_363_imag = _RAND_496[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_366_real = _RAND_497[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_366_imag = _RAND_498[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_369_real = _RAND_499[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_369_imag = _RAND_500[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_372_real = _RAND_501[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_372_imag = _RAND_502[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_375_real = _RAND_503[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_375_imag = _RAND_504[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_378_real = _RAND_505[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_378_imag = _RAND_506[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_381_real = _RAND_507[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_381_imag = _RAND_508[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_384_real = _RAND_509[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_384_imag = _RAND_510[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_387_real = _RAND_511[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_387_imag = _RAND_512[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_390_real = _RAND_513[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_390_imag = _RAND_514[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_393_real = _RAND_515[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_393_imag = _RAND_516[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_396_real = _RAND_517[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_396_imag = _RAND_518[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_399_real = _RAND_519[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_7__T_399_imag = _RAND_520[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_8_value = _RAND_521[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_sdf_stages_8__T_26 = _RAND_522[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_state = _RAND_523[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_initialOutDone = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_cnt = _RAND_525[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  fft_fft_SDFChainRadix22_cntValidOut = _RAND_526[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    fft_Queue__T_read[initvar] = _RAND_527[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_528 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    fft_Queue__T_data[initvar] = _RAND_528[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_529 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    fft_Queue__T_extra[initvar] = _RAND_529[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  fft_Queue_value = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  fft_Queue_value_1 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  fft_Queue__T_1 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  fft_busy = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    mag_logMagMux_magModule_Queue__T[initvar] = _RAND_534[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  mag_logMagMux_magModule_Queue_value = _RAND_535[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  mag_logMagMux_magModule_Queue_value_1 = _RAND_536[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  mag_logMagMux_magModule_Queue__T_1 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    mag_logMagMux_magModule_Queue_1__T[initvar] = _RAND_538[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  mag_logMagMux_magModule_Queue_1_value = _RAND_539[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  mag_logMagMux_magModule_Queue_1_value_1 = _RAND_540[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  mag_logMagMux_magModule_Queue_1__T_1 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_14 = _RAND_542[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  mag_logMagMux_magModule_jplMagOp1 = _RAND_543[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  mag_logMagMux_magModule_tmpOp2 = _RAND_544[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_18 = _RAND_545[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  mag_logMagMux_magModule_jplMagOp2 = _RAND_546[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_21 = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_24 = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  mag_logMagMux_magModule_squared_magnitude = _RAND_549[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_34 = _RAND_550[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_35 = _RAND_551[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  mag_logMagMux_magModule_queueCounter = _RAND_552[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_46 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_47 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_56 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_57 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  mag_logMagMux_magModule_queueCounter_1 = _RAND_557[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_64 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  mag_logMagMux_magModule__T_65 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    mag_Queue__T_read[initvar] = _RAND_560[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_561 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    mag_Queue__T_data[initvar] = _RAND_561[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_562 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    mag_Queue__T_extra[initvar] = _RAND_562[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  mag_Queue_value = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  mag_Queue_value_1 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  mag_Queue__T_1 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  mag_selReg = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    cfar_cfar_cfarCore_laggWindow_mem[initvar] = _RAND_567[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_568 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    cfar_cfar_cfarCore_laggWindow_outputQueue__T[initvar] = _RAND_568[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow_outputQueue__T_1 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow_writeIdxReg = _RAND_570[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow_last = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow_initialInDone = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow_validPrev = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_348 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_349 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_350 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_351 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_352 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_353 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_354 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_355 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_356 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_357 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_358 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_359 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_360 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_361 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_362 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_363 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_364 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_365 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_366 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_367 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_368 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_369 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_370 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_371 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_372 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_373 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_374 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_375 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_376 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_377 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_378 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_379 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_380 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_381 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_382 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_383 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_384 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_385 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_386 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_387 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_388 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_389 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_390 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_391 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_392 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_393 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_394 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_395 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_396 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_397 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_398 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_399 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_400 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_401 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_402 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_403 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_404 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_405 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_406 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_407 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_408 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_409 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_410 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_411 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggWindow__T_426 = _RAND_638[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_InitialInDone = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_last = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_0 = _RAND_641[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_1 = _RAND_642[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_2 = _RAND_643[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_3 = _RAND_644[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_4 = _RAND_645[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_5 = _RAND_646[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_6 = _RAND_647[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_7 = _RAND_648[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard_cntIn = _RAND_649[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_120 = _RAND_650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_121 = _RAND_651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_122 = _RAND_652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_123 = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_124 = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_125 = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_126 = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  cfar_cfar_cfarCore_laggGuard__T_127 = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  cfar_cfar_cfarCore_cellUnderTest_initialInDone = _RAND_658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  cfar_cfar_cfarCore_cellUnderTest_last = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  cfar_cfar_cfarCore_cellUnderTest_cut = _RAND_660[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  cfar_cfar_cfarCore_cellUnderTest_lastOut = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_InitialInDone = _RAND_662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_last = _RAND_663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_0 = _RAND_664[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_1 = _RAND_665[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_2 = _RAND_666[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_3 = _RAND_667[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_4 = _RAND_668[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_5 = _RAND_669[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_6 = _RAND_670[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_7 = _RAND_671[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard_cntIn = _RAND_672[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_120 = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_121 = _RAND_674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_122 = _RAND_675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_123 = _RAND_676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_124 = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_125 = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_126 = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadGuard__T_127 = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    cfar_cfar_cfarCore_leadWindow_mem[initvar] = _RAND_681[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_682 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    cfar_cfar_cfarCore_leadWindow_outputQueue__T[initvar] = _RAND_682[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow_outputQueue__T_1 = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow_writeIdxReg = _RAND_684[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow_last = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow_initialInDone = _RAND_686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow_validPrev = _RAND_687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_348 = _RAND_688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_349 = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_350 = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_351 = _RAND_691[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_352 = _RAND_692[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_353 = _RAND_693[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_354 = _RAND_694[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_355 = _RAND_695[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_356 = _RAND_696[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_357 = _RAND_697[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_358 = _RAND_698[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_359 = _RAND_699[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_360 = _RAND_700[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_361 = _RAND_701[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_362 = _RAND_702[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_363 = _RAND_703[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_364 = _RAND_704[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_365 = _RAND_705[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_366 = _RAND_706[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_367 = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_368 = _RAND_708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_369 = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_370 = _RAND_710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_371 = _RAND_711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_372 = _RAND_712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_373 = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_374 = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_375 = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_376 = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_377 = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_378 = _RAND_718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_379 = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_380 = _RAND_720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_381 = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_382 = _RAND_722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_383 = _RAND_723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_384 = _RAND_724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_385 = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_386 = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_387 = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_388 = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_389 = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_390 = _RAND_730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_391 = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_392 = _RAND_732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_393 = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_394 = _RAND_734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_395 = _RAND_735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_396 = _RAND_736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_397 = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_398 = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_399 = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_400 = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_401 = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_402 = _RAND_742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_403 = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_404 = _RAND_744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_405 = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_406 = _RAND_746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_407 = _RAND_747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_408 = _RAND_748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_409 = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_410 = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_411 = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leadWindow__T_426 = _RAND_752[15:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cfar_cfar_cfarCore_Queue__T_peak[initvar] = _RAND_753[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_754 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cfar_cfar_cfarCore_Queue__T_cut[initvar] = _RAND_754[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_755 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cfar_cfar_cfarCore_Queue__T_threshold[initvar] = _RAND_755[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  cfar_cfar_cfarCore_Queue_value = _RAND_756[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  cfar_cfar_cfarCore_Queue_value_1 = _RAND_757[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  cfar_cfar_cfarCore_Queue__T_1 = _RAND_758[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cfar_cfar_cfarCore_Queue_2__T[initvar] = _RAND_759[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  cfar_cfar_cfarCore_Queue_2_value = _RAND_760[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  cfar_cfar_cfarCore_Queue_2_value_1 = _RAND_761[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  cfar_cfar_cfarCore_Queue_2__T_1 = _RAND_762[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  cfar_cfar_cfarCore_lastCut = _RAND_763[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  cfar_cfar_cfarCore_flushing = _RAND_764[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  cfar_cfar_cfarCore_cntIn = _RAND_765[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  cfar_cfar_cfarCore_cntOut = _RAND_766[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  cfar_cfar_cfarCore_initialInDone = _RAND_767[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  cfar_cfar_cfarCore_sumlagg = _RAND_768[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  cfar_cfar_cfarCore_sumlead = _RAND_769[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  cfar_cfar_cfarCore_lastOut = _RAND_770[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  cfar_cfar_cfarCore_flushingDelayed = _RAND_771[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  cfar_cfar_cfarCore_enableRightThr = _RAND_772[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {2{`RANDOM}};
  cfar_cfar_cfarCore__T_94 = _RAND_773[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  cfar_cfar_cfarCore_cutDelayed = _RAND_774[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  cfar_cfar_cfarCore_leftNeighb = _RAND_775[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  cfar_cfar_cfarCore_rightNeighb = _RAND_776[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  cfar_cfar_cfarCore__T_106 = _RAND_777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  cfar_cfar_cfarCore__T_107 = _RAND_778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  cfar_cfar_cfarCore__T_120 = _RAND_779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  cfar_cfar_cfarCore__T_121 = _RAND_780[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cfar_Queue__T_read[initvar] = _RAND_781[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_782 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cfar_Queue__T_data[initvar] = _RAND_782[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_783 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cfar_Queue__T_extra[initvar] = _RAND_783[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  cfar_Queue_value = _RAND_784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  cfar_Queue_value_1 = _RAND_785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  cfar_Queue__T_1 = _RAND_786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  cfar_fftWin = _RAND_787[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  cfar_thresholdScaler = _RAND_788[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  cfar_peakGrouping = _RAND_789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  cfar_cfarMode = _RAND_790[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  cfar_windowCells = _RAND_791[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  cfar_guardCells = _RAND_792[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  cfar__T_6 = _RAND_793[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  widthAdapter_1__T_4 = _RAND_794[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  widthAdapter_1__T_10 = _RAND_795[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  widthAdapter_1__T_19 = _RAND_796[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  widthAdapter_1__T_26 = _RAND_797[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  widthAdapter_1__T_33 = _RAND_798[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_Queue__T_data[initvar] = _RAND_799[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_800 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_Queue__T_last[initvar] = _RAND_800[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  buffer_Queue_value = _RAND_801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  buffer_Queue_value_1 = _RAND_802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  buffer_Queue__T_1 = _RAND_803[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_1_Queue__T_data[initvar] = _RAND_804[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_805 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_1_Queue__T_last[initvar] = _RAND_805[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  buffer_1_Queue_value = _RAND_806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  buffer_1_Queue_value_1 = _RAND_807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  buffer_1_Queue__T_1 = _RAND_808[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_2_Queue__T_data[initvar] = _RAND_809[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_810 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_2_Queue__T_last[initvar] = _RAND_810[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  buffer_2_Queue_value = _RAND_811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  buffer_2_Queue_value_1 = _RAND_812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  buffer_2_Queue__T_1 = _RAND_813[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_814 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_3_Queue__T_data[initvar] = _RAND_814[47:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_815 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    buffer_3_Queue__T_last[initvar] = _RAND_815[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  buffer_3_Queue_value = _RAND_816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  buffer_3_Queue_value_1 = _RAND_817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  buffer_3_Queue__T_1 = _RAND_818[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    bus_awIn_0__T[initvar] = _RAND_819[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  bus_awIn_0_value = _RAND_820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  bus_awIn_0_value_1 = _RAND_821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  bus_awIn_0__T_1 = _RAND_822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  bus__T_59 = _RAND_823[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  bus__T_60 = _RAND_824[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  bus__T_302 = _RAND_825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  bus__T_373_0 = _RAND_826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  bus__T_373_1 = _RAND_827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  bus__T_373_2 = _RAND_828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  bus__T_313 = _RAND_829[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  bus__T_113 = _RAND_830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  bus__T_87 = _RAND_831[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  bus__T_88 = _RAND_832[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  bus__T_407 = _RAND_833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  bus__T_478_0 = _RAND_834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  bus__T_478_1 = _RAND_835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  bus__T_478_2 = _RAND_836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  bus__T_418 = _RAND_837[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge widthAdapter_clock) begin
    if (widthAdapter__T_10) begin
      widthAdapter__T <= widthAdapter_auto_in_bits_data;
    end
    if (widthAdapter__T_13) begin
      widthAdapter__T_1 <= widthAdapter_auto_in_bits_data;
    end
    if (widthAdapter__T_16) begin
      widthAdapter__T_2 <= widthAdapter_auto_in_bits_data;
    end
    if (widthAdapter_reset) begin
      widthAdapter__T_3 <= 2'h0;
    end else begin
      widthAdapter__T_3 <= widthAdapter__GEN_0[1:0];
    end
    if (widthAdapter__T_30) begin
      widthAdapter__T_20 <= widthAdapter_auto_in_bits_last;
    end
    if (widthAdapter__T_33) begin
      widthAdapter__T_21 <= widthAdapter_auto_in_bits_last;
    end
    if (widthAdapter__T_36) begin
      widthAdapter__T_22 <= widthAdapter_auto_in_bits_last;
    end
    if (widthAdapter_reset) begin
      widthAdapter__T_23 <= 2'h0;
    end else begin
      widthAdapter__T_23 <= widthAdapter__GEN_4[1:0];
    end
    if (widthAdapter_reset) begin
      widthAdapter__T_44 <= 2'h0;
    end else begin
      widthAdapter__T_44 <= widthAdapter__GEN_8[1:0];
    end
    if (widthAdapter_reset) begin
      widthAdapter__T_64 <= 2'h0;
    end else begin
      widthAdapter__T_64 <= widthAdapter__GEN_12[1:0];
    end
    if (widthAdapter_reset) begin
      widthAdapter__T_84 <= 2'h0;
    end else begin
      widthAdapter__T_84 <= widthAdapter__GEN_16[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter__T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter__T_104) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter__T_108) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter__T_108) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter__T_112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter__T_112) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter__T_116) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter__T_116) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_0_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_0_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_0_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_0_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_0_io_in_real;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_0_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_0_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_0_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_0_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_0_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_0_io_in_imag;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_0_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_0_butterfly_outputs_1_imag;
      end
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_1_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_1_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_1_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_1__T_21_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_1_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_1_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_1__T_21_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_1_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_1_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_1__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_1_io_in_real;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_1__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_1_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_1_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_1_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_1__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_1_io_in_imag;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_1__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_1_butterfly_outputs_1_imag;
      end
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_2_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_2_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_2__T_27_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_2_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_2__T_27_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_2_load_input) begin
        if (fft_fft_SDFChainRadix22__T_289) begin
          fft_fft_SDFChainRadix22_sdf_stages_2__T_21_real <= fft_fft_SDFChainRadix22_outputWires_1_imag;
        end else begin
          fft_fft_SDFChainRadix22_sdf_stages_2__T_21_real <= fft_fft_SDFChainRadix22_outputWires_1_real;
        end
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_2__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_2_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_2_load_input) begin
        if (fft_fft_SDFChainRadix22__T_289) begin
          fft_fft_SDFChainRadix22_sdf_stages_2__T_21_imag <= fft_fft_SDFChainRadix22__T_295;
        end else begin
          fft_fft_SDFChainRadix22_sdf_stages_2__T_21_imag <= fft_fft_SDFChainRadix22_outputWires_1_imag;
        end
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_2__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_2_butterfly_outputs_1_imag;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_2__T_24_real <= fft_fft_SDFChainRadix22_sdf_stages_2__T_21_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_2__T_24_imag <= fft_fft_SDFChainRadix22_sdf_stages_2__T_21_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_2__T_27_real <= fft_fft_SDFChainRadix22_sdf_stages_2__T_24_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_2_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_2__T_27_imag <= fft_fft_SDFChainRadix22_sdf_stages_2__T_24_imag;
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_3_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_3__T_39_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_3__T_39_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_3_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_3__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_3_io_in_real;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_3__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_3_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_3_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_3__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_3_io_in_imag;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_3__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_3_butterfly_outputs_1_imag;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_24_real <= fft_fft_SDFChainRadix22_sdf_stages_3__T_21_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_24_imag <= fft_fft_SDFChainRadix22_sdf_stages_3__T_21_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_27_real <= fft_fft_SDFChainRadix22_sdf_stages_3__T_24_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_27_imag <= fft_fft_SDFChainRadix22_sdf_stages_3__T_24_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_30_real <= fft_fft_SDFChainRadix22_sdf_stages_3__T_27_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_30_imag <= fft_fft_SDFChainRadix22_sdf_stages_3__T_27_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_33_real <= fft_fft_SDFChainRadix22_sdf_stages_3__T_30_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_33_imag <= fft_fft_SDFChainRadix22_sdf_stages_3__T_30_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_36_real <= fft_fft_SDFChainRadix22_sdf_stages_3__T_33_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_36_imag <= fft_fft_SDFChainRadix22_sdf_stages_3__T_33_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_39_real <= fft_fft_SDFChainRadix22_sdf_stages_3__T_36_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_3_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_3__T_39_imag <= fft_fft_SDFChainRadix22_sdf_stages_3__T_36_imag;
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_4_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_63_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_63_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_4_load_input) begin
        if (fft_fft_SDFChainRadix22__T_421) begin
          fft_fft_SDFChainRadix22_sdf_stages_4__T_21_real <= fft_fft_SDFChainRadix22_outputWires_3_imag;
        end else begin
          fft_fft_SDFChainRadix22_sdf_stages_4__T_21_real <= fft_fft_SDFChainRadix22_outputWires_3_real;
        end
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_4__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_4_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_4_load_input) begin
        if (fft_fft_SDFChainRadix22__T_421) begin
          fft_fft_SDFChainRadix22_sdf_stages_4__T_21_imag <= fft_fft_SDFChainRadix22__T_427;
        end else begin
          fft_fft_SDFChainRadix22_sdf_stages_4__T_21_imag <= fft_fft_SDFChainRadix22_outputWires_3_imag;
        end
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_4__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_4_butterfly_outputs_1_imag;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_24_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_21_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_24_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_21_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_27_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_24_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_27_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_24_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_30_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_27_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_30_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_27_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_33_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_30_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_33_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_30_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_36_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_33_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_36_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_33_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_39_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_36_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_39_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_36_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_42_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_39_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_42_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_39_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_45_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_42_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_45_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_42_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_48_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_45_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_48_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_45_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_51_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_48_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_51_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_48_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_54_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_51_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_54_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_51_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_57_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_54_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_57_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_54_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_60_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_57_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_60_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_57_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_63_real <= fft_fft_SDFChainRadix22_sdf_stages_4__T_60_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_4_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_4__T_63_imag <= fft_fft_SDFChainRadix22_sdf_stages_4__T_60_imag;
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_5_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_111_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_111_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_5_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_5__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_5_io_in_real;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_5__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_5_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_5_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_5__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_5_io_in_imag;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_5__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_5_butterfly_outputs_1_imag;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_24_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_21_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_24_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_21_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_27_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_24_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_27_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_24_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_30_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_27_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_30_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_27_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_33_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_30_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_33_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_30_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_36_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_33_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_36_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_33_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_39_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_36_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_39_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_36_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_42_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_39_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_42_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_39_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_45_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_42_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_45_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_42_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_48_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_45_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_48_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_45_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_51_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_48_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_51_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_48_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_54_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_51_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_54_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_51_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_57_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_54_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_57_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_54_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_60_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_57_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_60_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_57_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_63_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_60_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_63_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_60_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_66_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_63_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_66_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_63_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_69_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_66_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_69_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_66_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_72_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_69_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_72_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_69_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_75_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_72_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_75_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_72_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_78_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_75_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_78_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_75_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_81_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_78_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_81_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_78_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_84_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_81_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_84_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_81_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_87_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_84_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_87_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_84_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_90_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_87_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_90_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_87_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_93_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_90_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_93_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_90_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_96_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_93_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_96_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_93_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_99_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_96_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_99_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_96_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_102_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_99_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_102_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_99_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_105_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_102_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_105_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_102_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_108_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_105_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_108_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_105_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_111_real <= fft_fft_SDFChainRadix22_sdf_stages_5__T_108_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_5_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_5__T_111_imag <= fft_fft_SDFChainRadix22_sdf_stages_5__T_108_imag;
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_6_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_207_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_207_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_6_load_input) begin
        if (fft_fft_SDFChainRadix22__T_793) begin
          fft_fft_SDFChainRadix22_sdf_stages_6__T_21_real <= fft_fft_SDFChainRadix22_outputWires_5_imag;
        end else begin
          fft_fft_SDFChainRadix22_sdf_stages_6__T_21_real <= fft_fft_SDFChainRadix22_outputWires_5_real;
        end
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_6__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_6_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_6_load_input) begin
        if (fft_fft_SDFChainRadix22__T_793) begin
          fft_fft_SDFChainRadix22_sdf_stages_6__T_21_imag <= fft_fft_SDFChainRadix22__T_799;
        end else begin
          fft_fft_SDFChainRadix22_sdf_stages_6__T_21_imag <= fft_fft_SDFChainRadix22_outputWires_5_imag;
        end
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_6__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_6_butterfly_outputs_1_imag;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_24_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_21_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_24_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_21_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_27_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_24_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_27_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_24_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_30_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_27_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_30_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_27_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_33_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_30_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_33_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_30_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_36_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_33_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_36_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_33_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_39_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_36_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_39_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_36_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_42_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_39_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_42_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_39_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_45_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_42_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_45_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_42_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_48_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_45_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_48_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_45_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_51_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_48_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_51_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_48_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_54_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_51_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_54_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_51_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_57_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_54_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_57_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_54_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_60_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_57_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_60_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_57_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_63_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_60_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_63_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_60_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_66_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_63_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_66_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_63_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_69_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_66_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_69_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_66_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_72_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_69_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_72_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_69_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_75_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_72_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_75_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_72_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_78_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_75_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_78_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_75_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_81_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_78_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_81_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_78_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_84_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_81_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_84_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_81_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_87_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_84_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_87_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_84_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_90_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_87_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_90_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_87_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_93_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_90_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_93_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_90_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_96_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_93_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_96_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_93_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_99_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_96_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_99_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_96_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_102_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_99_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_102_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_99_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_105_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_102_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_105_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_102_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_108_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_105_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_108_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_105_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_111_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_108_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_111_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_108_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_114_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_111_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_114_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_111_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_117_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_114_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_117_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_114_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_120_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_117_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_120_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_117_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_123_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_120_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_123_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_120_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_126_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_123_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_126_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_123_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_129_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_126_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_129_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_126_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_132_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_129_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_132_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_129_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_135_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_132_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_135_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_132_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_138_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_135_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_138_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_135_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_141_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_138_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_141_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_138_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_144_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_141_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_144_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_141_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_147_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_144_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_147_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_144_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_150_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_147_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_150_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_147_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_153_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_150_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_153_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_150_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_156_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_153_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_156_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_153_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_159_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_156_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_159_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_156_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_162_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_159_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_162_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_159_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_165_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_162_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_165_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_162_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_168_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_165_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_168_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_165_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_171_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_168_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_171_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_168_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_174_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_171_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_174_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_171_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_177_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_174_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_177_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_174_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_180_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_177_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_180_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_177_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_183_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_180_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_183_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_180_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_186_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_183_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_186_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_183_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_189_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_186_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_189_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_186_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_192_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_189_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_192_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_189_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_195_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_192_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_195_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_192_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_198_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_195_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_198_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_195_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_201_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_198_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_201_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_198_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_204_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_201_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_204_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_201_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_207_real <= fft_fft_SDFChainRadix22_sdf_stages_6__T_204_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_6_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_6__T_207_imag <= fft_fft_SDFChainRadix22_sdf_stages_6__T_204_imag;
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_7_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7_feedback_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_399_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7_feedback_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_399_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_7_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_7__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_7_io_in_real;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_7__T_21_real <= fft_fft_SDFChainRadix22_sdf_stages_7_butterfly_outputs_1_real;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      if (fft_fft_SDFChainRadix22_sdf_stages_7_load_input) begin
        fft_fft_SDFChainRadix22_sdf_stages_7__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_7_io_in_imag;
      end else begin
        fft_fft_SDFChainRadix22_sdf_stages_7__T_21_imag <= fft_fft_SDFChainRadix22_sdf_stages_7_butterfly_outputs_1_imag;
      end
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_24_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_21_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_24_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_21_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_27_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_24_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_27_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_24_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_30_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_27_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_30_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_27_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_33_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_30_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_33_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_30_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_36_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_33_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_36_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_33_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_39_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_36_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_39_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_36_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_42_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_39_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_42_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_39_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_45_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_42_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_45_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_42_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_48_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_45_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_48_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_45_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_51_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_48_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_51_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_48_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_54_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_51_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_54_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_51_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_57_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_54_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_57_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_54_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_60_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_57_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_60_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_57_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_63_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_60_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_63_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_60_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_66_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_63_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_66_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_63_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_69_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_66_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_69_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_66_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_72_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_69_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_72_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_69_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_75_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_72_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_75_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_72_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_78_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_75_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_78_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_75_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_81_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_78_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_81_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_78_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_84_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_81_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_84_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_81_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_87_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_84_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_87_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_84_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_90_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_87_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_90_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_87_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_93_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_90_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_93_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_90_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_96_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_93_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_96_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_93_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_99_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_96_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_99_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_96_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_102_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_99_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_102_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_99_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_105_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_102_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_105_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_102_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_108_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_105_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_108_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_105_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_111_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_108_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_111_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_108_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_114_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_111_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_114_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_111_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_117_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_114_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_117_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_114_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_120_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_117_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_120_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_117_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_123_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_120_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_123_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_120_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_126_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_123_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_126_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_123_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_129_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_126_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_129_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_126_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_132_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_129_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_132_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_129_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_135_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_132_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_135_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_132_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_138_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_135_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_138_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_135_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_141_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_138_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_141_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_138_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_144_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_141_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_144_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_141_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_147_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_144_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_147_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_144_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_150_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_147_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_150_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_147_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_153_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_150_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_153_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_150_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_156_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_153_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_156_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_153_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_159_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_156_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_159_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_156_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_162_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_159_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_162_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_159_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_165_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_162_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_165_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_162_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_168_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_165_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_168_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_165_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_171_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_168_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_171_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_168_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_174_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_171_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_174_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_171_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_177_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_174_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_177_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_174_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_180_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_177_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_180_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_177_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_183_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_180_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_183_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_180_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_186_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_183_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_186_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_183_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_189_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_186_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_189_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_186_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_192_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_189_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_192_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_189_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_195_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_192_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_195_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_192_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_198_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_195_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_198_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_195_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_201_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_198_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_201_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_198_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_204_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_201_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_204_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_201_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_207_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_204_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_207_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_204_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_210_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_207_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_210_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_207_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_213_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_210_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_213_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_210_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_216_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_213_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_216_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_213_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_219_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_216_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_219_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_216_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_222_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_219_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_222_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_219_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_225_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_222_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_225_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_222_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_228_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_225_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_228_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_225_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_231_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_228_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_231_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_228_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_234_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_231_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_234_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_231_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_237_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_234_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_237_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_234_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_240_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_237_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_240_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_237_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_243_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_240_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_243_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_240_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_246_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_243_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_246_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_243_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_249_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_246_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_249_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_246_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_252_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_249_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_252_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_249_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_255_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_252_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_255_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_252_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_258_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_255_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_258_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_255_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_261_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_258_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_261_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_258_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_264_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_261_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_264_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_261_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_267_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_264_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_267_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_264_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_270_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_267_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_270_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_267_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_273_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_270_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_273_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_270_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_276_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_273_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_276_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_273_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_279_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_276_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_279_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_276_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_282_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_279_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_282_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_279_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_285_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_282_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_285_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_282_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_288_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_285_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_288_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_285_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_291_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_288_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_291_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_288_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_294_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_291_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_294_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_291_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_297_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_294_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_297_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_294_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_300_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_297_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_300_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_297_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_303_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_300_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_303_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_300_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_306_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_303_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_306_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_303_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_309_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_306_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_309_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_306_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_312_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_309_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_312_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_309_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_315_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_312_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_315_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_312_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_318_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_315_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_318_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_315_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_321_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_318_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_321_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_318_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_324_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_321_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_324_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_321_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_327_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_324_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_327_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_324_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_330_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_327_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_330_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_327_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_333_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_330_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_333_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_330_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_336_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_333_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_336_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_333_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_339_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_336_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_339_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_336_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_342_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_339_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_342_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_339_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_345_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_342_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_345_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_342_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_348_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_345_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_348_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_345_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_351_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_348_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_351_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_348_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_354_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_351_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_354_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_351_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_357_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_354_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_357_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_354_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_360_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_357_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_360_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_357_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_363_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_360_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_363_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_360_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_366_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_363_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_366_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_363_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_369_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_366_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_369_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_366_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_372_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_369_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_372_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_369_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_375_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_372_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_375_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_372_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_378_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_375_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_378_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_375_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_381_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_378_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_381_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_378_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_384_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_381_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_384_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_381_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_387_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_384_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_387_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_384_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_390_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_387_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_390_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_387_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_393_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_390_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_393_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_390_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_396_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_393_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_396_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_393_imag;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_399_real <= fft_fft_SDFChainRadix22_sdf_stages_7__T_396_real;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_7_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_7__T_399_imag <= fft_fft_SDFChainRadix22_sdf_stages_7__T_396_imag;
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_sdf_stages_8_clock) begin
    if (fft_fft_SDFChainRadix22_sdf_stages_8_reset) begin
      fft_fft_SDFChainRadix22_sdf_stages_8_value <= 8'h0;
    end else if (fft_fft_SDFChainRadix22_sdf_stages_8_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_8_value <= fft_fft_SDFChainRadix22_sdf_stages_8__T_22;
    end
    if (fft_fft_SDFChainRadix22_sdf_stages_8_reset) begin
      fft_fft_SDFChainRadix22_sdf_stages_8__T_26 <= 8'hff;
    end else if (fft_fft_SDFChainRadix22_sdf_stages_8_io_en) begin
      fft_fft_SDFChainRadix22_sdf_stages_8__T_26 <= fft_fft_SDFChainRadix22_sdf_stages_8_value;
    end
  end
  always @(posedge fft_fft_SDFChainRadix22_clock) begin
    if (fft_fft_SDFChainRadix22_reset) begin
      fft_fft_SDFChainRadix22_state <= 2'h0;
    end else if (fft_fft_SDFChainRadix22__T_53) begin
      if (fft_fft_SDFChainRadix22__T_46) begin
        fft_fft_SDFChainRadix22_state <= 2'h1;
      end
    end else if (fft_fft_SDFChainRadix22__T_56) begin
      if (fft_fft_SDFChainRadix22_fireLast) begin
        fft_fft_SDFChainRadix22_state <= 2'h2;
      end
    end else if (fft_fft_SDFChainRadix22__T_57) begin
      if (fft_fft_SDFChainRadix22_io_lastOut) begin
        fft_fft_SDFChainRadix22_state <= 2'h0;
      end
    end
    if (fft_fft_SDFChainRadix22_reset) begin
      fft_fft_SDFChainRadix22_initialOutDone <= 1'h0;
    end else begin
      fft_fft_SDFChainRadix22_initialOutDone <= fft_fft_SDFChainRadix22__GEN_46;
    end
    if (fft_fft_SDFChainRadix22_reset) begin
      fft_fft_SDFChainRadix22_cnt <= 10'h0;
    end else if (fft_fft_SDFChainRadix22__T_62) begin
      fft_fft_SDFChainRadix22_cnt <= 10'h0;
    end else if (fft_fft_SDFChainRadix22_enableInit) begin
      fft_fft_SDFChainRadix22_cnt <= fft_fft_SDFChainRadix22__T_125;
    end
    if (fft_fft_SDFChainRadix22_reset) begin
      fft_fft_SDFChainRadix22_cntValidOut <= 9'h0;
    end else if (fft_fft_SDFChainRadix22__T_77) begin
      fft_fft_SDFChainRadix22_cntValidOut <= 9'h0;
    end else if (fft_fft_SDFChainRadix22__T_61) begin
      fft_fft_SDFChainRadix22_cntValidOut <= fft_fft_SDFChainRadix22__T_80;
    end
  end
  always @(posedge fft_Queue_clock) begin
    if(fft_Queue__T_read__T_10_en & fft_Queue__T_read__T_10_mask) begin
      fft_Queue__T_read[fft_Queue__T_read__T_10_addr] <= fft_Queue__T_read__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(fft_Queue__T_data__T_10_en & fft_Queue__T_data__T_10_mask) begin
      fft_Queue__T_data[fft_Queue__T_data__T_10_addr] <= fft_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(fft_Queue__T_extra__T_10_en & fft_Queue__T_extra__T_10_mask) begin
      fft_Queue__T_extra[fft_Queue__T_extra__T_10_addr] <= fft_Queue__T_extra__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (fft_Queue_reset) begin
      fft_Queue_value <= 1'h0;
    end else if (fft_Queue__T_6) begin
      fft_Queue_value <= fft_Queue__T_12;
    end
    if (fft_Queue_reset) begin
      fft_Queue_value_1 <= 1'h0;
    end else if (fft_Queue__T_8) begin
      fft_Queue_value_1 <= fft_Queue__T_14;
    end
    if (fft_Queue_reset) begin
      fft_Queue__T_1 <= 1'h0;
    end else if (fft_Queue__T_15) begin
      fft_Queue__T_1 <= fft_Queue__T_6;
    end
  end
  always @(posedge fft_clock) begin
    if (fft_reset) begin
      fft_busy <= 1'h0;
    end else begin
      fft_busy <= fft_fft_io_busy;
    end
  end
  always @(posedge mag_logMagMux_magModule_Queue_clock) begin
    if(mag_logMagMux_magModule_Queue__T__T_10_en & mag_logMagMux_magModule_Queue__T__T_10_mask) begin
      mag_logMagMux_magModule_Queue__T[mag_logMagMux_magModule_Queue__T__T_10_addr] <= mag_logMagMux_magModule_Queue__T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (mag_logMagMux_magModule_Queue_reset) begin
      mag_logMagMux_magModule_Queue_value <= 2'h0;
    end else if (mag_logMagMux_magModule_Queue__T_6) begin
      mag_logMagMux_magModule_Queue_value <= mag_logMagMux_magModule_Queue__T_12;
    end
    if (mag_logMagMux_magModule_Queue_reset) begin
      mag_logMagMux_magModule_Queue_value_1 <= 2'h0;
    end else if (mag_logMagMux_magModule_Queue__T_8) begin
      mag_logMagMux_magModule_Queue_value_1 <= mag_logMagMux_magModule_Queue__T_14;
    end
    if (mag_logMagMux_magModule_Queue_reset) begin
      mag_logMagMux_magModule_Queue__T_1 <= 1'h0;
    end else if (mag_logMagMux_magModule_Queue__T_15) begin
      mag_logMagMux_magModule_Queue__T_1 <= mag_logMagMux_magModule_Queue__T_6;
    end
  end
  always @(posedge mag_logMagMux_magModule_Queue_1_clock) begin
    if(mag_logMagMux_magModule_Queue_1__T__T_10_en & mag_logMagMux_magModule_Queue_1__T__T_10_mask) begin
      mag_logMagMux_magModule_Queue_1__T[mag_logMagMux_magModule_Queue_1__T__T_10_addr] <= mag_logMagMux_magModule_Queue_1__T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (mag_logMagMux_magModule_Queue_1_reset) begin
      mag_logMagMux_magModule_Queue_1_value <= 2'h0;
    end else if (mag_logMagMux_magModule_Queue_1__T_6) begin
      mag_logMagMux_magModule_Queue_1_value <= mag_logMagMux_magModule_Queue_1__T_12;
    end
    if (mag_logMagMux_magModule_Queue_1_reset) begin
      mag_logMagMux_magModule_Queue_1_value_1 <= 2'h0;
    end else if (mag_logMagMux_magModule_Queue_1__T_8) begin
      mag_logMagMux_magModule_Queue_1_value_1 <= mag_logMagMux_magModule_Queue_1__T_14;
    end
    if (mag_logMagMux_magModule_Queue_1_reset) begin
      mag_logMagMux_magModule_Queue_1__T_1 <= 1'h0;
    end else if (mag_logMagMux_magModule_Queue_1__T_15) begin
      mag_logMagMux_magModule_Queue_1__T_1 <= mag_logMagMux_magModule_Queue_1__T_6;
    end
  end
  always @(posedge mag_logMagMux_magModule_clock) begin
    mag_logMagMux_magModule__T_14 <= $signed(mag_logMagMux_magModule_u) + $signed(mag_logMagMux_magModule__GEN_16);
    mag_logMagMux_magModule_jplMagOp1 <= mag_logMagMux_magModule__T_14;
    mag_logMagMux_magModule_tmpOp2 <= $signed(mag_logMagMux_magModule_u) - $signed(mag_logMagMux_magModule__GEN_17);
    mag_logMagMux_magModule__T_18 <= mag_logMagMux_magModule_v[15:1];
    mag_logMagMux_magModule_jplMagOp2 <= $signed(mag_logMagMux_magModule_tmpOp2) + $signed(mag_logMagMux_magModule__GEN_18);
    mag_logMagMux_magModule__T_21 <= $signed(mag_logMagMux_magModule_absInReal) * $signed(mag_logMagMux_magModule_absInReal);
    mag_logMagMux_magModule__T_24 <= $signed(mag_logMagMux_magModule_absInImag) * $signed(mag_logMagMux_magModule_absInImag);
    mag_logMagMux_magModule_squared_magnitude <= $signed(mag_logMagMux_magModule__T_22) + $signed(mag_logMagMux_magModule__T_25);
    mag_logMagMux_magModule__T_34 <= mag_logMagMux_magModule_io_sel;
    mag_logMagMux_magModule__T_35 <= mag_logMagMux_magModule__T_34;
    if (mag_logMagMux_magModule_reset) begin
      mag_logMagMux_magModule_queueCounter <= 2'h0;
    end else begin
      mag_logMagMux_magModule_queueCounter <= mag_logMagMux_magModule__T_43[1:0];
    end
    if (mag_logMagMux_magModule_reset) begin
      mag_logMagMux_magModule__T_46 <= 1'h0;
    end else begin
      mag_logMagMux_magModule__T_46 <= mag_logMagMux_magModule__T_40;
    end
    if (mag_logMagMux_magModule_reset) begin
      mag_logMagMux_magModule__T_47 <= 1'h0;
    end else begin
      mag_logMagMux_magModule__T_47 <= mag_logMagMux_magModule__T_46;
    end
    mag_logMagMux_magModule__T_56 <= mag_logMagMux_magModule_io_lastIn & mag_logMagMux_magModule__T_54;
    mag_logMagMux_magModule__T_57 <= mag_logMagMux_magModule__T_56;
    if (mag_logMagMux_magModule_reset) begin
      mag_logMagMux_magModule_queueCounter_1 <= 2'h0;
    end else begin
      mag_logMagMux_magModule_queueCounter_1 <= mag_logMagMux_magModule__T_61[1:0];
    end
    if (mag_logMagMux_magModule_reset) begin
      mag_logMagMux_magModule__T_64 <= 1'h0;
    end else begin
      mag_logMagMux_magModule__T_64 <= mag_logMagMux_magModule__T_58;
    end
    if (mag_logMagMux_magModule_reset) begin
      mag_logMagMux_magModule__T_65 <= 1'h0;
    end else begin
      mag_logMagMux_magModule__T_65 <= mag_logMagMux_magModule__T_64;
    end
  end
  always @(posedge mag_Queue_clock) begin
    if(mag_Queue__T_read__T_10_en & mag_Queue__T_read__T_10_mask) begin
      mag_Queue__T_read[mag_Queue__T_read__T_10_addr] <= mag_Queue__T_read__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(mag_Queue__T_data__T_10_en & mag_Queue__T_data__T_10_mask) begin
      mag_Queue__T_data[mag_Queue__T_data__T_10_addr] <= mag_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(mag_Queue__T_extra__T_10_en & mag_Queue__T_extra__T_10_mask) begin
      mag_Queue__T_extra[mag_Queue__T_extra__T_10_addr] <= mag_Queue__T_extra__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (mag_Queue_reset) begin
      mag_Queue_value <= 1'h0;
    end else if (mag_Queue__T_6) begin
      mag_Queue_value <= mag_Queue__T_12;
    end
    if (mag_Queue_reset) begin
      mag_Queue_value_1 <= 1'h0;
    end else if (mag_Queue__T_8) begin
      mag_Queue_value_1 <= mag_Queue__T_14;
    end
    if (mag_Queue_reset) begin
      mag_Queue__T_1 <= 1'h0;
    end else if (mag_Queue__T_15) begin
      mag_Queue__T_1 <= mag_Queue__T_6;
    end
  end
  always @(posedge mag_clock) begin
    if (mag_reset) begin
      mag_selReg <= 1'h0;
    end else if (mag__T_98) begin
      mag_selReg <= mag__T_100;
    end
  end
  always @(posedge cfar_cfar_cfarCore_laggWindow_clock) begin
    if(cfar_cfar_cfarCore_laggWindow_mem__T_418_en & cfar_cfar_cfarCore_laggWindow_mem__T_418_mask) begin
      cfar_cfar_cfarCore_laggWindow_mem[cfar_cfar_cfarCore_laggWindow_mem__T_418_addr] <= cfar_cfar_cfarCore_laggWindow_mem__T_418_data; // @[CFARUtils.scala 505:26]
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow_writeIdxReg <= 6'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_417) begin
      if (cfar_cfar_cfarCore_laggWindow__T_419) begin
        cfar_cfar_cfarCore_laggWindow_writeIdxReg <= cfar_cfar_cfarCore_laggWindow__T_3;
      end else begin
        cfar_cfar_cfarCore_laggWindow_writeIdxReg <= 6'h0;
      end
    end else if (cfar_cfar_cfarCore_laggWindow_resetAll) begin
      cfar_cfar_cfarCore_laggWindow_writeIdxReg <= 6'h0;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow_last <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow_resetAll) begin
      cfar_cfar_cfarCore_laggWindow_last <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_laggWindow_last <= cfar_cfar_cfarCore_laggWindow__GEN_2;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow_initialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow_resetAll) begin
      cfar_cfar_cfarCore_laggWindow_initialInDone <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_laggWindow_initialInDone <= cfar_cfar_cfarCore_laggWindow__GEN_1;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow_validPrev <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_laggWindow_validPrev <= cfar_cfar_cfarCore_laggWindow_io_in_valid;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_348 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_21) begin
      cfar_cfar_cfarCore_laggWindow__T_348 <= cfar_cfar_cfarCore_laggWindow_fireLastIn;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_349 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_346) begin
      cfar_cfar_cfarCore_laggWindow__T_349 <= cfar_cfar_cfarCore_laggWindow__T_348;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_350 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_345) begin
      cfar_cfar_cfarCore_laggWindow__T_350 <= cfar_cfar_cfarCore_laggWindow__T_349;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_351 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_344) begin
      cfar_cfar_cfarCore_laggWindow__T_351 <= cfar_cfar_cfarCore_laggWindow__T_350;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_352 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_343) begin
      cfar_cfar_cfarCore_laggWindow__T_352 <= cfar_cfar_cfarCore_laggWindow__T_351;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_353 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_342) begin
      cfar_cfar_cfarCore_laggWindow__T_353 <= cfar_cfar_cfarCore_laggWindow__T_352;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_354 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_341) begin
      cfar_cfar_cfarCore_laggWindow__T_354 <= cfar_cfar_cfarCore_laggWindow__T_353;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_355 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_340) begin
      cfar_cfar_cfarCore_laggWindow__T_355 <= cfar_cfar_cfarCore_laggWindow__T_354;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_356 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_339) begin
      cfar_cfar_cfarCore_laggWindow__T_356 <= cfar_cfar_cfarCore_laggWindow__T_355;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_357 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_338) begin
      cfar_cfar_cfarCore_laggWindow__T_357 <= cfar_cfar_cfarCore_laggWindow__T_356;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_358 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_337) begin
      cfar_cfar_cfarCore_laggWindow__T_358 <= cfar_cfar_cfarCore_laggWindow__T_357;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_359 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_336) begin
      cfar_cfar_cfarCore_laggWindow__T_359 <= cfar_cfar_cfarCore_laggWindow__T_358;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_360 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_335) begin
      cfar_cfar_cfarCore_laggWindow__T_360 <= cfar_cfar_cfarCore_laggWindow__T_359;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_361 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_334) begin
      cfar_cfar_cfarCore_laggWindow__T_361 <= cfar_cfar_cfarCore_laggWindow__T_360;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_362 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_333) begin
      cfar_cfar_cfarCore_laggWindow__T_362 <= cfar_cfar_cfarCore_laggWindow__T_361;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_363 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_332) begin
      cfar_cfar_cfarCore_laggWindow__T_363 <= cfar_cfar_cfarCore_laggWindow__T_362;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_364 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_331) begin
      cfar_cfar_cfarCore_laggWindow__T_364 <= cfar_cfar_cfarCore_laggWindow__T_363;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_365 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_330) begin
      cfar_cfar_cfarCore_laggWindow__T_365 <= cfar_cfar_cfarCore_laggWindow__T_364;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_366 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_329) begin
      cfar_cfar_cfarCore_laggWindow__T_366 <= cfar_cfar_cfarCore_laggWindow__T_365;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_367 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_328) begin
      cfar_cfar_cfarCore_laggWindow__T_367 <= cfar_cfar_cfarCore_laggWindow__T_366;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_368 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_327) begin
      cfar_cfar_cfarCore_laggWindow__T_368 <= cfar_cfar_cfarCore_laggWindow__T_367;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_369 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_326) begin
      cfar_cfar_cfarCore_laggWindow__T_369 <= cfar_cfar_cfarCore_laggWindow__T_368;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_370 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_325) begin
      cfar_cfar_cfarCore_laggWindow__T_370 <= cfar_cfar_cfarCore_laggWindow__T_369;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_371 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_324) begin
      cfar_cfar_cfarCore_laggWindow__T_371 <= cfar_cfar_cfarCore_laggWindow__T_370;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_372 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_323) begin
      cfar_cfar_cfarCore_laggWindow__T_372 <= cfar_cfar_cfarCore_laggWindow__T_371;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_373 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_322) begin
      cfar_cfar_cfarCore_laggWindow__T_373 <= cfar_cfar_cfarCore_laggWindow__T_372;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_374 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_321) begin
      cfar_cfar_cfarCore_laggWindow__T_374 <= cfar_cfar_cfarCore_laggWindow__T_373;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_375 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_320) begin
      cfar_cfar_cfarCore_laggWindow__T_375 <= cfar_cfar_cfarCore_laggWindow__T_374;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_376 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_319) begin
      cfar_cfar_cfarCore_laggWindow__T_376 <= cfar_cfar_cfarCore_laggWindow__T_375;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_377 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_318) begin
      cfar_cfar_cfarCore_laggWindow__T_377 <= cfar_cfar_cfarCore_laggWindow__T_376;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_378 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_317) begin
      cfar_cfar_cfarCore_laggWindow__T_378 <= cfar_cfar_cfarCore_laggWindow__T_377;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_379 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_316) begin
      cfar_cfar_cfarCore_laggWindow__T_379 <= cfar_cfar_cfarCore_laggWindow__T_378;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_380 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_315) begin
      cfar_cfar_cfarCore_laggWindow__T_380 <= cfar_cfar_cfarCore_laggWindow__T_379;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_381 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_314) begin
      cfar_cfar_cfarCore_laggWindow__T_381 <= cfar_cfar_cfarCore_laggWindow__T_380;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_382 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_313) begin
      cfar_cfar_cfarCore_laggWindow__T_382 <= cfar_cfar_cfarCore_laggWindow__T_381;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_383 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_312) begin
      cfar_cfar_cfarCore_laggWindow__T_383 <= cfar_cfar_cfarCore_laggWindow__T_382;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_384 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_311) begin
      cfar_cfar_cfarCore_laggWindow__T_384 <= cfar_cfar_cfarCore_laggWindow__T_383;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_385 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_310) begin
      cfar_cfar_cfarCore_laggWindow__T_385 <= cfar_cfar_cfarCore_laggWindow__T_384;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_386 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_309) begin
      cfar_cfar_cfarCore_laggWindow__T_386 <= cfar_cfar_cfarCore_laggWindow__T_385;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_387 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_308) begin
      cfar_cfar_cfarCore_laggWindow__T_387 <= cfar_cfar_cfarCore_laggWindow__T_386;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_388 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_307) begin
      cfar_cfar_cfarCore_laggWindow__T_388 <= cfar_cfar_cfarCore_laggWindow__T_387;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_389 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_306) begin
      cfar_cfar_cfarCore_laggWindow__T_389 <= cfar_cfar_cfarCore_laggWindow__T_388;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_390 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_305) begin
      cfar_cfar_cfarCore_laggWindow__T_390 <= cfar_cfar_cfarCore_laggWindow__T_389;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_391 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_304) begin
      cfar_cfar_cfarCore_laggWindow__T_391 <= cfar_cfar_cfarCore_laggWindow__T_390;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_392 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_303) begin
      cfar_cfar_cfarCore_laggWindow__T_392 <= cfar_cfar_cfarCore_laggWindow__T_391;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_393 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_302) begin
      cfar_cfar_cfarCore_laggWindow__T_393 <= cfar_cfar_cfarCore_laggWindow__T_392;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_394 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_301) begin
      cfar_cfar_cfarCore_laggWindow__T_394 <= cfar_cfar_cfarCore_laggWindow__T_393;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_395 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_300) begin
      cfar_cfar_cfarCore_laggWindow__T_395 <= cfar_cfar_cfarCore_laggWindow__T_394;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_396 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_299) begin
      cfar_cfar_cfarCore_laggWindow__T_396 <= cfar_cfar_cfarCore_laggWindow__T_395;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_397 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_298) begin
      cfar_cfar_cfarCore_laggWindow__T_397 <= cfar_cfar_cfarCore_laggWindow__T_396;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_398 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_297) begin
      cfar_cfar_cfarCore_laggWindow__T_398 <= cfar_cfar_cfarCore_laggWindow__T_397;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_399 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_296) begin
      cfar_cfar_cfarCore_laggWindow__T_399 <= cfar_cfar_cfarCore_laggWindow__T_398;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_400 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_295) begin
      cfar_cfar_cfarCore_laggWindow__T_400 <= cfar_cfar_cfarCore_laggWindow__T_399;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_401 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_294) begin
      cfar_cfar_cfarCore_laggWindow__T_401 <= cfar_cfar_cfarCore_laggWindow__T_400;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_402 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_293) begin
      cfar_cfar_cfarCore_laggWindow__T_402 <= cfar_cfar_cfarCore_laggWindow__T_401;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_403 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_292) begin
      cfar_cfar_cfarCore_laggWindow__T_403 <= cfar_cfar_cfarCore_laggWindow__T_402;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_404 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_291) begin
      cfar_cfar_cfarCore_laggWindow__T_404 <= cfar_cfar_cfarCore_laggWindow__T_403;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_405 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_290) begin
      cfar_cfar_cfarCore_laggWindow__T_405 <= cfar_cfar_cfarCore_laggWindow__T_404;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_406 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_289) begin
      cfar_cfar_cfarCore_laggWindow__T_406 <= cfar_cfar_cfarCore_laggWindow__T_405;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_407 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_288) begin
      cfar_cfar_cfarCore_laggWindow__T_407 <= cfar_cfar_cfarCore_laggWindow__T_406;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_408 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_287) begin
      cfar_cfar_cfarCore_laggWindow__T_408 <= cfar_cfar_cfarCore_laggWindow__T_407;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_409 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_286) begin
      cfar_cfar_cfarCore_laggWindow__T_409 <= cfar_cfar_cfarCore_laggWindow__T_408;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_410 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_285) begin
      cfar_cfar_cfarCore_laggWindow__T_410 <= cfar_cfar_cfarCore_laggWindow__T_409;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_411 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow__T_284) begin
      cfar_cfar_cfarCore_laggWindow__T_411 <= cfar_cfar_cfarCore_laggWindow__T_410;
    end
    if (cfar_cfar_cfarCore_laggWindow_reset) begin
      cfar_cfar_cfarCore_laggWindow__T_426 <= 16'sh0;
    end else begin
      cfar_cfar_cfarCore_laggWindow__T_426 <= cfar_cfar_cfarCore_laggWindow_mem__T_423_data;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore_laggWindow__T_25) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:330 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 330:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore_laggWindow__T_25) begin
          $fatal; // @[CFARUtils.scala 330:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge cfar_cfar_cfarCore_laggWindow_outputQueue_clock) begin
    if(cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_en & cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_mask) begin
      cfar_cfar_cfarCore_laggWindow_outputQueue__T[cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_addr] <= cfar_cfar_cfarCore_laggWindow_outputQueue__T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (cfar_cfar_cfarCore_laggWindow_outputQueue_reset) begin
      cfar_cfar_cfarCore_laggWindow_outputQueue__T_1 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggWindow_outputQueue__T_11) begin
      if (cfar_cfar_cfarCore_laggWindow_outputQueue__T_3) begin
        if (cfar_cfar_cfarCore_laggWindow_outputQueue_io_deq_ready) begin
          cfar_cfar_cfarCore_laggWindow_outputQueue__T_1 <= 1'h0;
        end else begin
          cfar_cfar_cfarCore_laggWindow_outputQueue__T_1 <= cfar_cfar_cfarCore_laggWindow_outputQueue__T_6;
        end
      end else begin
        cfar_cfar_cfarCore_laggWindow_outputQueue__T_1 <= cfar_cfar_cfarCore_laggWindow_outputQueue__T_6;
      end
    end
  end
  always @(posedge cfar_cfar_cfarCore_laggGuard_clock) begin
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_InitialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_132) begin
      cfar_cfar_cfarCore_laggGuard_InitialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_63) begin
      cfar_cfar_cfarCore_laggGuard_InitialInDone <= cfar_cfar_cfarCore_laggGuard__GEN_10;
    end else begin
      cfar_cfar_cfarCore_laggGuard_InitialInDone <= cfar_cfar_cfarCore_laggGuard__GEN_11;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_last <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_132) begin
      cfar_cfar_cfarCore_laggGuard_last <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_laggGuard_last <= cfar_cfar_cfarCore_laggGuard__GEN_8;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_0 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_46) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_0 <= cfar_cfar_cfarCore_laggGuard_io_in_bits;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_1 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_45) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_1 <= cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_0;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_2 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_44) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_2 <= cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_1;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_3 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_43) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_3 <= cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_2;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_4 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_42) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_4 <= cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_3;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_5 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_41) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_5 <= cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_4;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_6 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_40) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_6 <= cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_5;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_7 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_39) begin
      cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_7 <= cfar_cfar_cfarCore_laggGuard_adjShiftRegOut_6;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard_cntIn <= 4'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_132) begin
      cfar_cfar_cfarCore_laggGuard_cntIn <= 4'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_1) begin
      cfar_cfar_cfarCore_laggGuard_cntIn <= cfar_cfar_cfarCore_laggGuard__T_62;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_120 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_73) begin
      cfar_cfar_cfarCore_laggGuard__T_120 <= cfar_cfar_cfarCore_laggGuard__T_59;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_121 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_118) begin
      cfar_cfar_cfarCore_laggGuard__T_121 <= cfar_cfar_cfarCore_laggGuard__T_120;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_122 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_117) begin
      cfar_cfar_cfarCore_laggGuard__T_122 <= cfar_cfar_cfarCore_laggGuard__T_121;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_123 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_116) begin
      cfar_cfar_cfarCore_laggGuard__T_123 <= cfar_cfar_cfarCore_laggGuard__T_122;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_124 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_115) begin
      cfar_cfar_cfarCore_laggGuard__T_124 <= cfar_cfar_cfarCore_laggGuard__T_123;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_125 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_114) begin
      cfar_cfar_cfarCore_laggGuard__T_125 <= cfar_cfar_cfarCore_laggGuard__T_124;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_126 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_113) begin
      cfar_cfar_cfarCore_laggGuard__T_126 <= cfar_cfar_cfarCore_laggGuard__T_125;
    end
    if (cfar_cfar_cfarCore_laggGuard_reset) begin
      cfar_cfar_cfarCore_laggGuard__T_127 <= 1'h0;
    end else if (cfar_cfar_cfarCore_laggGuard__T_112) begin
      cfar_cfar_cfarCore_laggGuard__T_127 <= cfar_cfar_cfarCore_laggGuard__T_126;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore_laggGuard__T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:345 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 345:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore_laggGuard__T_6) begin
          $fatal; // @[CFARUtils.scala 345:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore_laggGuard__T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:330 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 330:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore_laggGuard__T_6) begin
          $fatal; // @[CFARUtils.scala 330:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge cfar_cfar_cfarCore_cellUnderTest_clock) begin
    if (cfar_cfar_cfarCore_cellUnderTest_reset) begin
      cfar_cfar_cfarCore_cellUnderTest_initialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_cellUnderTest__T_9) begin
      cfar_cfar_cfarCore_cellUnderTest_initialInDone <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_cellUnderTest_initialInDone <= cfar_cfar_cfarCore_cellUnderTest__GEN_0;
    end
    if (cfar_cfar_cfarCore_cellUnderTest_reset) begin
      cfar_cfar_cfarCore_cellUnderTest_last <= 1'h0;
    end else if (cfar_cfar_cfarCore_cellUnderTest__T_9) begin
      cfar_cfar_cfarCore_cellUnderTest_last <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_cellUnderTest_last <= cfar_cfar_cfarCore_cellUnderTest__GEN_2;
    end
    if (cfar_cfar_cfarCore_cellUnderTest_reset) begin
      cfar_cfar_cfarCore_cellUnderTest_cut <= 16'sh0;
    end else if (cfar_cfar_cfarCore_cellUnderTest_en) begin
      cfar_cfar_cfarCore_cellUnderTest_cut <= cfar_cfar_cfarCore_cellUnderTest_io_in_bits;
    end
    if (cfar_cfar_cfarCore_cellUnderTest_reset) begin
      cfar_cfar_cfarCore_cellUnderTest_lastOut <= 1'h0;
    end else if (cfar_cfar_cfarCore_cellUnderTest_io_out_ready) begin
      cfar_cfar_cfarCore_cellUnderTest_lastOut <= cfar_cfar_cfarCore_cellUnderTest__T_7;
    end
  end
  always @(posedge cfar_cfar_cfarCore_leadGuard_clock) begin
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_InitialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_132) begin
      cfar_cfar_cfarCore_leadGuard_InitialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_63) begin
      cfar_cfar_cfarCore_leadGuard_InitialInDone <= cfar_cfar_cfarCore_leadGuard__GEN_10;
    end else begin
      cfar_cfar_cfarCore_leadGuard_InitialInDone <= cfar_cfar_cfarCore_leadGuard__GEN_11;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_last <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_132) begin
      cfar_cfar_cfarCore_leadGuard_last <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_leadGuard_last <= cfar_cfar_cfarCore_leadGuard__GEN_8;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_0 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_46) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_0 <= cfar_cfar_cfarCore_leadGuard_io_in_bits;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_1 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_45) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_1 <= cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_0;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_2 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_44) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_2 <= cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_1;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_3 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_43) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_3 <= cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_2;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_4 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_42) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_4 <= cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_3;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_5 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_41) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_5 <= cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_4;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_6 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_40) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_6 <= cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_5;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_7 <= 16'sh0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_39) begin
      cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_7 <= cfar_cfar_cfarCore_leadGuard_adjShiftRegOut_6;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard_cntIn <= 4'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_132) begin
      cfar_cfar_cfarCore_leadGuard_cntIn <= 4'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_1) begin
      cfar_cfar_cfarCore_leadGuard_cntIn <= cfar_cfar_cfarCore_leadGuard__T_62;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_120 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_73) begin
      cfar_cfar_cfarCore_leadGuard__T_120 <= cfar_cfar_cfarCore_leadGuard__T_59;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_121 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_118) begin
      cfar_cfar_cfarCore_leadGuard__T_121 <= cfar_cfar_cfarCore_leadGuard__T_120;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_122 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_117) begin
      cfar_cfar_cfarCore_leadGuard__T_122 <= cfar_cfar_cfarCore_leadGuard__T_121;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_123 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_116) begin
      cfar_cfar_cfarCore_leadGuard__T_123 <= cfar_cfar_cfarCore_leadGuard__T_122;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_124 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_115) begin
      cfar_cfar_cfarCore_leadGuard__T_124 <= cfar_cfar_cfarCore_leadGuard__T_123;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_125 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_114) begin
      cfar_cfar_cfarCore_leadGuard__T_125 <= cfar_cfar_cfarCore_leadGuard__T_124;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_126 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_113) begin
      cfar_cfar_cfarCore_leadGuard__T_126 <= cfar_cfar_cfarCore_leadGuard__T_125;
    end
    if (cfar_cfar_cfarCore_leadGuard_reset) begin
      cfar_cfar_cfarCore_leadGuard__T_127 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadGuard__T_112) begin
      cfar_cfar_cfarCore_leadGuard__T_127 <= cfar_cfar_cfarCore_leadGuard__T_126;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore_leadGuard__T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:345 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 345:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore_leadGuard__T_6) begin
          $fatal; // @[CFARUtils.scala 345:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore_leadGuard__T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:330 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 330:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore_leadGuard__T_6) begin
          $fatal; // @[CFARUtils.scala 330:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge cfar_cfar_cfarCore_leadWindow_clock) begin
    if(cfar_cfar_cfarCore_leadWindow_mem__T_418_en & cfar_cfar_cfarCore_leadWindow_mem__T_418_mask) begin
      cfar_cfar_cfarCore_leadWindow_mem[cfar_cfar_cfarCore_leadWindow_mem__T_418_addr] <= cfar_cfar_cfarCore_leadWindow_mem__T_418_data; // @[CFARUtils.scala 505:26]
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow_writeIdxReg <= 6'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_417) begin
      if (cfar_cfar_cfarCore_leadWindow__T_419) begin
        cfar_cfar_cfarCore_leadWindow_writeIdxReg <= cfar_cfar_cfarCore_leadWindow__T_3;
      end else begin
        cfar_cfar_cfarCore_leadWindow_writeIdxReg <= 6'h0;
      end
    end else if (cfar_cfar_cfarCore_leadWindow_resetAll) begin
      cfar_cfar_cfarCore_leadWindow_writeIdxReg <= 6'h0;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow_last <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow_resetAll) begin
      cfar_cfar_cfarCore_leadWindow_last <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_leadWindow_last <= cfar_cfar_cfarCore_leadWindow__GEN_2;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow_initialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow_resetAll) begin
      cfar_cfar_cfarCore_leadWindow_initialInDone <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_leadWindow_initialInDone <= cfar_cfar_cfarCore_leadWindow__GEN_1;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow_validPrev <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_leadWindow_validPrev <= cfar_cfar_cfarCore_leadWindow_io_in_valid;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_348 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_21) begin
      cfar_cfar_cfarCore_leadWindow__T_348 <= cfar_cfar_cfarCore_leadWindow_fireLastIn;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_349 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_346) begin
      cfar_cfar_cfarCore_leadWindow__T_349 <= cfar_cfar_cfarCore_leadWindow__T_348;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_350 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_345) begin
      cfar_cfar_cfarCore_leadWindow__T_350 <= cfar_cfar_cfarCore_leadWindow__T_349;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_351 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_344) begin
      cfar_cfar_cfarCore_leadWindow__T_351 <= cfar_cfar_cfarCore_leadWindow__T_350;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_352 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_343) begin
      cfar_cfar_cfarCore_leadWindow__T_352 <= cfar_cfar_cfarCore_leadWindow__T_351;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_353 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_342) begin
      cfar_cfar_cfarCore_leadWindow__T_353 <= cfar_cfar_cfarCore_leadWindow__T_352;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_354 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_341) begin
      cfar_cfar_cfarCore_leadWindow__T_354 <= cfar_cfar_cfarCore_leadWindow__T_353;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_355 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_340) begin
      cfar_cfar_cfarCore_leadWindow__T_355 <= cfar_cfar_cfarCore_leadWindow__T_354;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_356 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_339) begin
      cfar_cfar_cfarCore_leadWindow__T_356 <= cfar_cfar_cfarCore_leadWindow__T_355;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_357 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_338) begin
      cfar_cfar_cfarCore_leadWindow__T_357 <= cfar_cfar_cfarCore_leadWindow__T_356;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_358 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_337) begin
      cfar_cfar_cfarCore_leadWindow__T_358 <= cfar_cfar_cfarCore_leadWindow__T_357;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_359 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_336) begin
      cfar_cfar_cfarCore_leadWindow__T_359 <= cfar_cfar_cfarCore_leadWindow__T_358;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_360 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_335) begin
      cfar_cfar_cfarCore_leadWindow__T_360 <= cfar_cfar_cfarCore_leadWindow__T_359;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_361 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_334) begin
      cfar_cfar_cfarCore_leadWindow__T_361 <= cfar_cfar_cfarCore_leadWindow__T_360;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_362 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_333) begin
      cfar_cfar_cfarCore_leadWindow__T_362 <= cfar_cfar_cfarCore_leadWindow__T_361;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_363 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_332) begin
      cfar_cfar_cfarCore_leadWindow__T_363 <= cfar_cfar_cfarCore_leadWindow__T_362;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_364 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_331) begin
      cfar_cfar_cfarCore_leadWindow__T_364 <= cfar_cfar_cfarCore_leadWindow__T_363;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_365 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_330) begin
      cfar_cfar_cfarCore_leadWindow__T_365 <= cfar_cfar_cfarCore_leadWindow__T_364;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_366 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_329) begin
      cfar_cfar_cfarCore_leadWindow__T_366 <= cfar_cfar_cfarCore_leadWindow__T_365;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_367 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_328) begin
      cfar_cfar_cfarCore_leadWindow__T_367 <= cfar_cfar_cfarCore_leadWindow__T_366;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_368 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_327) begin
      cfar_cfar_cfarCore_leadWindow__T_368 <= cfar_cfar_cfarCore_leadWindow__T_367;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_369 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_326) begin
      cfar_cfar_cfarCore_leadWindow__T_369 <= cfar_cfar_cfarCore_leadWindow__T_368;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_370 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_325) begin
      cfar_cfar_cfarCore_leadWindow__T_370 <= cfar_cfar_cfarCore_leadWindow__T_369;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_371 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_324) begin
      cfar_cfar_cfarCore_leadWindow__T_371 <= cfar_cfar_cfarCore_leadWindow__T_370;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_372 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_323) begin
      cfar_cfar_cfarCore_leadWindow__T_372 <= cfar_cfar_cfarCore_leadWindow__T_371;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_373 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_322) begin
      cfar_cfar_cfarCore_leadWindow__T_373 <= cfar_cfar_cfarCore_leadWindow__T_372;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_374 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_321) begin
      cfar_cfar_cfarCore_leadWindow__T_374 <= cfar_cfar_cfarCore_leadWindow__T_373;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_375 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_320) begin
      cfar_cfar_cfarCore_leadWindow__T_375 <= cfar_cfar_cfarCore_leadWindow__T_374;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_376 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_319) begin
      cfar_cfar_cfarCore_leadWindow__T_376 <= cfar_cfar_cfarCore_leadWindow__T_375;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_377 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_318) begin
      cfar_cfar_cfarCore_leadWindow__T_377 <= cfar_cfar_cfarCore_leadWindow__T_376;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_378 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_317) begin
      cfar_cfar_cfarCore_leadWindow__T_378 <= cfar_cfar_cfarCore_leadWindow__T_377;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_379 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_316) begin
      cfar_cfar_cfarCore_leadWindow__T_379 <= cfar_cfar_cfarCore_leadWindow__T_378;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_380 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_315) begin
      cfar_cfar_cfarCore_leadWindow__T_380 <= cfar_cfar_cfarCore_leadWindow__T_379;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_381 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_314) begin
      cfar_cfar_cfarCore_leadWindow__T_381 <= cfar_cfar_cfarCore_leadWindow__T_380;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_382 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_313) begin
      cfar_cfar_cfarCore_leadWindow__T_382 <= cfar_cfar_cfarCore_leadWindow__T_381;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_383 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_312) begin
      cfar_cfar_cfarCore_leadWindow__T_383 <= cfar_cfar_cfarCore_leadWindow__T_382;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_384 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_311) begin
      cfar_cfar_cfarCore_leadWindow__T_384 <= cfar_cfar_cfarCore_leadWindow__T_383;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_385 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_310) begin
      cfar_cfar_cfarCore_leadWindow__T_385 <= cfar_cfar_cfarCore_leadWindow__T_384;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_386 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_309) begin
      cfar_cfar_cfarCore_leadWindow__T_386 <= cfar_cfar_cfarCore_leadWindow__T_385;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_387 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_308) begin
      cfar_cfar_cfarCore_leadWindow__T_387 <= cfar_cfar_cfarCore_leadWindow__T_386;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_388 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_307) begin
      cfar_cfar_cfarCore_leadWindow__T_388 <= cfar_cfar_cfarCore_leadWindow__T_387;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_389 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_306) begin
      cfar_cfar_cfarCore_leadWindow__T_389 <= cfar_cfar_cfarCore_leadWindow__T_388;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_390 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_305) begin
      cfar_cfar_cfarCore_leadWindow__T_390 <= cfar_cfar_cfarCore_leadWindow__T_389;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_391 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_304) begin
      cfar_cfar_cfarCore_leadWindow__T_391 <= cfar_cfar_cfarCore_leadWindow__T_390;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_392 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_303) begin
      cfar_cfar_cfarCore_leadWindow__T_392 <= cfar_cfar_cfarCore_leadWindow__T_391;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_393 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_302) begin
      cfar_cfar_cfarCore_leadWindow__T_393 <= cfar_cfar_cfarCore_leadWindow__T_392;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_394 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_301) begin
      cfar_cfar_cfarCore_leadWindow__T_394 <= cfar_cfar_cfarCore_leadWindow__T_393;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_395 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_300) begin
      cfar_cfar_cfarCore_leadWindow__T_395 <= cfar_cfar_cfarCore_leadWindow__T_394;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_396 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_299) begin
      cfar_cfar_cfarCore_leadWindow__T_396 <= cfar_cfar_cfarCore_leadWindow__T_395;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_397 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_298) begin
      cfar_cfar_cfarCore_leadWindow__T_397 <= cfar_cfar_cfarCore_leadWindow__T_396;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_398 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_297) begin
      cfar_cfar_cfarCore_leadWindow__T_398 <= cfar_cfar_cfarCore_leadWindow__T_397;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_399 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_296) begin
      cfar_cfar_cfarCore_leadWindow__T_399 <= cfar_cfar_cfarCore_leadWindow__T_398;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_400 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_295) begin
      cfar_cfar_cfarCore_leadWindow__T_400 <= cfar_cfar_cfarCore_leadWindow__T_399;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_401 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_294) begin
      cfar_cfar_cfarCore_leadWindow__T_401 <= cfar_cfar_cfarCore_leadWindow__T_400;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_402 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_293) begin
      cfar_cfar_cfarCore_leadWindow__T_402 <= cfar_cfar_cfarCore_leadWindow__T_401;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_403 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_292) begin
      cfar_cfar_cfarCore_leadWindow__T_403 <= cfar_cfar_cfarCore_leadWindow__T_402;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_404 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_291) begin
      cfar_cfar_cfarCore_leadWindow__T_404 <= cfar_cfar_cfarCore_leadWindow__T_403;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_405 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_290) begin
      cfar_cfar_cfarCore_leadWindow__T_405 <= cfar_cfar_cfarCore_leadWindow__T_404;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_406 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_289) begin
      cfar_cfar_cfarCore_leadWindow__T_406 <= cfar_cfar_cfarCore_leadWindow__T_405;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_407 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_288) begin
      cfar_cfar_cfarCore_leadWindow__T_407 <= cfar_cfar_cfarCore_leadWindow__T_406;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_408 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_287) begin
      cfar_cfar_cfarCore_leadWindow__T_408 <= cfar_cfar_cfarCore_leadWindow__T_407;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_409 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_286) begin
      cfar_cfar_cfarCore_leadWindow__T_409 <= cfar_cfar_cfarCore_leadWindow__T_408;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_410 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_285) begin
      cfar_cfar_cfarCore_leadWindow__T_410 <= cfar_cfar_cfarCore_leadWindow__T_409;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_411 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow__T_284) begin
      cfar_cfar_cfarCore_leadWindow__T_411 <= cfar_cfar_cfarCore_leadWindow__T_410;
    end
    if (cfar_cfar_cfarCore_leadWindow_reset) begin
      cfar_cfar_cfarCore_leadWindow__T_426 <= 16'sh0;
    end else begin
      cfar_cfar_cfarCore_leadWindow__T_426 <= cfar_cfar_cfarCore_leadWindow_mem__T_423_data;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore_leadWindow__T_25) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:330 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 330:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore_leadWindow__T_25) begin
          $fatal; // @[CFARUtils.scala 330:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge cfar_cfar_cfarCore_leadWindow_outputQueue_clock) begin
    if(cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_en & cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_mask) begin
      cfar_cfar_cfarCore_leadWindow_outputQueue__T[cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_addr] <= cfar_cfar_cfarCore_leadWindow_outputQueue__T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (cfar_cfar_cfarCore_leadWindow_outputQueue_reset) begin
      cfar_cfar_cfarCore_leadWindow_outputQueue__T_1 <= 1'h0;
    end else if (cfar_cfar_cfarCore_leadWindow_outputQueue__T_11) begin
      if (cfar_cfar_cfarCore_leadWindow_outputQueue__T_3) begin
        if (cfar_cfar_cfarCore_leadWindow_outputQueue_io_deq_ready) begin
          cfar_cfar_cfarCore_leadWindow_outputQueue__T_1 <= 1'h0;
        end else begin
          cfar_cfar_cfarCore_leadWindow_outputQueue__T_1 <= cfar_cfar_cfarCore_leadWindow_outputQueue__T_6;
        end
      end else begin
        cfar_cfar_cfarCore_leadWindow_outputQueue__T_1 <= cfar_cfar_cfarCore_leadWindow_outputQueue__T_6;
      end
    end
  end
  always @(posedge cfar_cfar_cfarCore_Queue_clock) begin
    if(cfar_cfar_cfarCore_Queue__T_peak__T_10_en & cfar_cfar_cfarCore_Queue__T_peak__T_10_mask) begin
      cfar_cfar_cfarCore_Queue__T_peak[cfar_cfar_cfarCore_Queue__T_peak__T_10_addr] <= cfar_cfar_cfarCore_Queue__T_peak__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(cfar_cfar_cfarCore_Queue__T_cut__T_10_en & cfar_cfar_cfarCore_Queue__T_cut__T_10_mask) begin
      cfar_cfar_cfarCore_Queue__T_cut[cfar_cfar_cfarCore_Queue__T_cut__T_10_addr] <= cfar_cfar_cfarCore_Queue__T_cut__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(cfar_cfar_cfarCore_Queue__T_threshold__T_10_en & cfar_cfar_cfarCore_Queue__T_threshold__T_10_mask) begin
      cfar_cfar_cfarCore_Queue__T_threshold[cfar_cfar_cfarCore_Queue__T_threshold__T_10_addr] <= cfar_cfar_cfarCore_Queue__T_threshold__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (cfar_cfar_cfarCore_Queue_reset) begin
      cfar_cfar_cfarCore_Queue_value <= 1'h0;
    end else if (cfar_cfar_cfarCore_Queue__GEN_16) begin
      cfar_cfar_cfarCore_Queue_value <= cfar_cfar_cfarCore_Queue__T_12;
    end
    if (cfar_cfar_cfarCore_Queue_reset) begin
      cfar_cfar_cfarCore_Queue_value_1 <= 1'h0;
    end else if (cfar_cfar_cfarCore_Queue__GEN_15) begin
      cfar_cfar_cfarCore_Queue_value_1 <= cfar_cfar_cfarCore_Queue__T_14;
    end
    if (cfar_cfar_cfarCore_Queue_reset) begin
      cfar_cfar_cfarCore_Queue__T_1 <= 1'h0;
    end else if (cfar_cfar_cfarCore_Queue__T_15) begin
      if (cfar_cfar_cfarCore_Queue__T_4) begin
        if (cfar_cfar_cfarCore_Queue_io_deq_ready) begin
          cfar_cfar_cfarCore_Queue__T_1 <= 1'h0;
        end else begin
          cfar_cfar_cfarCore_Queue__T_1 <= cfar_cfar_cfarCore_Queue__T_6;
        end
      end else begin
        cfar_cfar_cfarCore_Queue__T_1 <= cfar_cfar_cfarCore_Queue__T_6;
      end
    end
  end
  always @(posedge cfar_cfar_cfarCore_Queue_2_clock) begin
    if(cfar_cfar_cfarCore_Queue_2__T__T_10_en & cfar_cfar_cfarCore_Queue_2__T__T_10_mask) begin
      cfar_cfar_cfarCore_Queue_2__T[cfar_cfar_cfarCore_Queue_2__T__T_10_addr] <= cfar_cfar_cfarCore_Queue_2__T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (cfar_cfar_cfarCore_Queue_2_reset) begin
      cfar_cfar_cfarCore_Queue_2_value <= 1'h0;
    end else if (cfar_cfar_cfarCore_Queue_2__GEN_12) begin
      cfar_cfar_cfarCore_Queue_2_value <= cfar_cfar_cfarCore_Queue_2__T_12;
    end
    if (cfar_cfar_cfarCore_Queue_2_reset) begin
      cfar_cfar_cfarCore_Queue_2_value_1 <= 1'h0;
    end else if (cfar_cfar_cfarCore_Queue_2__GEN_11) begin
      cfar_cfar_cfarCore_Queue_2_value_1 <= cfar_cfar_cfarCore_Queue_2__T_14;
    end
    if (cfar_cfar_cfarCore_Queue_2_reset) begin
      cfar_cfar_cfarCore_Queue_2__T_1 <= 1'h0;
    end else if (cfar_cfar_cfarCore_Queue_2__T_15) begin
      if (cfar_cfar_cfarCore_Queue_2__T_4) begin
        if (cfar_cfar_cfarCore_Queue_2_io_deq_ready) begin
          cfar_cfar_cfarCore_Queue_2__T_1 <= 1'h0;
        end else begin
          cfar_cfar_cfarCore_Queue_2__T_1 <= cfar_cfar_cfarCore_Queue_2__T_6;
        end
      end else begin
        cfar_cfar_cfarCore_Queue_2__T_1 <= cfar_cfar_cfarCore_Queue_2__T_6;
      end
    end
  end
  always @(posedge cfar_cfar_cfarCore_clock) begin
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_lastCut <= 1'h0;
    end else if (cfar_cfar_cfarCore__T_43) begin
      cfar_cfar_cfarCore_lastCut <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_lastCut <= cfar_cfar_cfarCore__GEN_9;
    end
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_flushing <= 1'h0;
    end else if (cfar_cfar_cfarCore_io_lastOut) begin
      cfar_cfar_cfarCore_flushing <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_flushing <= cfar_cfar_cfarCore__GEN_6;
    end
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_cntIn <= 9'h0;
    end else if (cfar_cfar_cfarCore__T_30) begin
      cfar_cfar_cfarCore_cntIn <= 9'h0;
    end else if (cfar_cfar_cfarCore__T_21) begin
      cfar_cfar_cfarCore_cntIn <= cfar_cfar_cfarCore__T_23;
    end
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_cntOut <= 9'h0;
    end else if (cfar_cfar_cfarCore__T_41) begin
      cfar_cfar_cfarCore_cntOut <= 9'h0;
    end else if (cfar_cfar_cfarCore__T_29) begin
      cfar_cfar_cfarCore_cntOut <= cfar_cfar_cfarCore__T_33;
    end
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_initialInDone <= 1'h0;
    end else if (cfar_cfar_cfarCore_io_lastOut) begin
      cfar_cfar_cfarCore_initialInDone <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_initialInDone <= cfar_cfar_cfarCore__GEN_2;
    end
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_sumlagg <= 20'sh0;
    end else if (cfar_cfar_cfarCore_io_lastOut) begin
      cfar_cfar_cfarCore_sumlagg <= 20'sh0;
    end else if (cfar_cfar_cfarCore__T_21) begin
      if (cfar_cfar_cfarCore_laggWindow_io_memFull) begin
        if (cfar_cfar_cfarCore__T_47) begin
          cfar_cfar_cfarCore_sumlagg <= cfar_cfar_cfarCore__T_53;
        end
      end else begin
        cfar_cfar_cfarCore_sumlagg <= cfar_cfar_cfarCore__T_50;
      end
    end
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_sumlead <= 20'sh0;
    end else if (cfar_cfar_cfarCore_lastCut) begin
      cfar_cfar_cfarCore_sumlead <= 20'sh0;
    end else if (cfar_cfar_cfarCore__T_59) begin
      if (cfar_cfar_cfarCore_leadWindow_io_memFull) begin
        if (cfar_cfar_cfarCore__T_60) begin
          cfar_cfar_cfarCore_sumlead <= cfar_cfar_cfarCore__T_66;
        end
      end else begin
        cfar_cfar_cfarCore_sumlead <= cfar_cfar_cfarCore__T_63;
      end
    end
    cfar_cfar_cfarCore_lastOut <= cfar_cfar_cfarCore_cellUnderTest_io_lastOut;
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_flushingDelayed <= 1'h0;
    end else if (cfar_cfar_cfarCore_io_lastOut) begin
      cfar_cfar_cfarCore_flushingDelayed <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_flushingDelayed <= cfar_cfar_cfarCore_flushing;
    end
    if (cfar_cfar_cfarCore_reset) begin
      cfar_cfar_cfarCore_enableRightThr <= 1'h0;
    end else if (cfar_cfar_cfarCore_io_lastOut) begin
      cfar_cfar_cfarCore_enableRightThr <= 1'h0;
    end else begin
      cfar_cfar_cfarCore_enableRightThr <= cfar_cfar_cfarCore__GEN_21;
    end
    cfar_cfar_cfarCore__T_94 <= $signed(cfar_cfar_cfarCore_thrWithoutScaling) * $signed(cfar_cfar_cfarCore__GEN_51);
    cfar_cfar_cfarCore_cutDelayed <= cfar_cfar_cfarCore_cellUnderTest_io_out_bits;
    if (3'h7 == cfar_cfar_cfarCore__T_97) begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_7;
    end else if (3'h6 == cfar_cfar_cfarCore__T_97) begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_6;
    end else if (3'h5 == cfar_cfar_cfarCore__T_97) begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_5;
    end else if (3'h4 == cfar_cfar_cfarCore__T_97) begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_4;
    end else if (3'h3 == cfar_cfar_cfarCore__T_97) begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_3;
    end else if (3'h2 == cfar_cfar_cfarCore__T_97) begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_2;
    end else if (3'h1 == cfar_cfar_cfarCore__T_97) begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_1;
    end else begin
      cfar_cfar_cfarCore_leftNeighb <= cfar_cfar_cfarCore__GEN_25;
    end
    cfar_cfar_cfarCore_rightNeighb <= cfar_cfar_cfarCore_laggGuard_io_parallelOut_0;
    cfar_cfar_cfarCore__T_106 <= cfar_cfar_cfarCore_initialInDone & cfar_cfar_cfarCore__T_21;
    cfar_cfar_cfarCore__T_107 <= cfar_cfar_cfarCore_io_out_ready;
    cfar_cfar_cfarCore__T_120 <= cfar_cfar_cfarCore_initialInDone & cfar_cfar_cfarCore__T_21;
    cfar_cfar_cfarCore__T_121 <= cfar_cfar_cfarCore_io_out_ready;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore__T_10) begin
          $fwrite(32'h80000002,"Assertion failed: FFT size must be larger than total number of shifting cells inside CFAR core\n    at CFARCoreWithMem.scala:33 assert(io.fftWin > 2.U * io.windowCells + 2.U * io.guardCells + 1.U, \"FFT size must be larger than total number of shifting cells inside CFAR core\")\n"); // @[CFARCoreWithMem.scala 33:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore__T_10) begin
          $fatal; // @[CFARCoreWithMem.scala 33:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (cfar_cfar_cfarCore__T_14) begin
          $fwrite(32'h80000002,"Assertion failed: Number of guard cells should be greater than 0\n    at CFARCoreWithMem.scala:34 assert(io.guardCells > 0.U, \"Number of guard cells should be greater than 0\")\n"); // @[CFARCoreWithMem.scala 34:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (cfar_cfar_cfarCore__T_14) begin
          $fatal; // @[CFARCoreWithMem.scala 34:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge cfar_Queue_clock) begin
    if(cfar_Queue__T_read__T_10_en & cfar_Queue__T_read__T_10_mask) begin
      cfar_Queue__T_read[cfar_Queue__T_read__T_10_addr] <= cfar_Queue__T_read__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(cfar_Queue__T_data__T_10_en & cfar_Queue__T_data__T_10_mask) begin
      cfar_Queue__T_data[cfar_Queue__T_data__T_10_addr] <= cfar_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(cfar_Queue__T_extra__T_10_en & cfar_Queue__T_extra__T_10_mask) begin
      cfar_Queue__T_extra[cfar_Queue__T_extra__T_10_addr] <= cfar_Queue__T_extra__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (cfar_Queue_reset) begin
      cfar_Queue_value <= 1'h0;
    end else if (cfar_Queue__T_6) begin
      cfar_Queue_value <= cfar_Queue__T_12;
    end
    if (cfar_Queue_reset) begin
      cfar_Queue_value_1 <= 1'h0;
    end else if (cfar_Queue__T_8) begin
      cfar_Queue_value_1 <= cfar_Queue__T_14;
    end
    if (cfar_Queue_reset) begin
      cfar_Queue__T_1 <= 1'h0;
    end else if (cfar_Queue__T_15) begin
      cfar_Queue__T_1 <= cfar_Queue__T_6;
    end
  end
  always @(posedge cfar_clock) begin
    if (cfar_reset) begin
      cfar_fftWin <= 10'h200;
    end else if (cfar__T_121) begin
      cfar_fftWin <= cfar__T_123;
    end
    if (cfar_reset) begin
      cfar_thresholdScaler <= 16'h0;
    end else if (cfar__T_167) begin
      cfar_thresholdScaler <= cfar__T_169;
    end
    if (cfar_reset) begin
      cfar_peakGrouping <= 1'h0;
    end else if (cfar__T_213) begin
      cfar_peakGrouping <= cfar__T_215;
    end
    if (cfar_reset) begin
      cfar_cfarMode <= 2'h0;
    end else if (cfar__T_236) begin
      cfar_cfarMode <= cfar__T_238;
    end
    if (cfar_reset) begin
      cfar_windowCells <= 7'h40;
    end else if (cfar__T_259) begin
      cfar_windowCells <= cfar__T_261;
    end
    if (cfar_reset) begin
      cfar_guardCells <= 4'h8;
    end else if (cfar__T_144) begin
      cfar_guardCells <= cfar__T_146;
    end
    if (cfar_reset) begin
      cfar__T_6 <= 3'h0;
    end else if (cfar__T_190) begin
      cfar__T_6 <= cfar__T_192;
    end
  end
  always @(posedge widthAdapter_1_clock) begin
    if (widthAdapter_1_reset) begin
      widthAdapter_1__T_4 <= 2'h0;
    end else begin
      widthAdapter_1__T_4 <= widthAdapter_1__GEN_0[1:0];
    end
    if (widthAdapter_1_reset) begin
      widthAdapter_1__T_10 <= 2'h0;
    end else begin
      widthAdapter_1__T_10 <= widthAdapter_1__GEN_1[1:0];
    end
    if (widthAdapter_1_reset) begin
      widthAdapter_1__T_19 <= 2'h0;
    end else begin
      widthAdapter_1__T_19 <= widthAdapter_1__GEN_2[1:0];
    end
    if (widthAdapter_1_reset) begin
      widthAdapter_1__T_26 <= 2'h0;
    end else begin
      widthAdapter_1__T_26 <= widthAdapter_1__GEN_3[1:0];
    end
    if (widthAdapter_1_reset) begin
      widthAdapter_1__T_33 <= 2'h0;
    end else begin
      widthAdapter_1__T_33 <= widthAdapter_1__GEN_4[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter_1__T_58) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:46 assert(ir0 === ir1)\n"); // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter_1__T_58) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter_1__T_62) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:47 assert(ir0 === ir2)\n"); // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter_1__T_62) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter_1__T_66) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:48 assert(ir0 === ir3)\n"); // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter_1__T_66) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (widthAdapter_1__T_70) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:49 assert(ir0 === ir4)\n"); // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (widthAdapter_1__T_70) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge buffer_Queue_clock) begin
    if(buffer_Queue__T_data__T_10_en & buffer_Queue__T_data__T_10_mask) begin
      buffer_Queue__T_data[buffer_Queue__T_data__T_10_addr] <= buffer_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(buffer_Queue__T_last__T_10_en & buffer_Queue__T_last__T_10_mask) begin
      buffer_Queue__T_last[buffer_Queue__T_last__T_10_addr] <= buffer_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (buffer_Queue_reset) begin
      buffer_Queue_value <= 1'h0;
    end else if (buffer_Queue__T_6) begin
      buffer_Queue_value <= buffer_Queue__T_12;
    end
    if (buffer_Queue_reset) begin
      buffer_Queue_value_1 <= 1'h0;
    end else if (buffer_Queue__T_8) begin
      buffer_Queue_value_1 <= buffer_Queue__T_14;
    end
    if (buffer_Queue_reset) begin
      buffer_Queue__T_1 <= 1'h0;
    end else if (buffer_Queue__T_15) begin
      buffer_Queue__T_1 <= buffer_Queue__T_6;
    end
  end
  always @(posedge buffer_1_Queue_clock) begin
    if(buffer_1_Queue__T_data__T_10_en & buffer_1_Queue__T_data__T_10_mask) begin
      buffer_1_Queue__T_data[buffer_1_Queue__T_data__T_10_addr] <= buffer_1_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(buffer_1_Queue__T_last__T_10_en & buffer_1_Queue__T_last__T_10_mask) begin
      buffer_1_Queue__T_last[buffer_1_Queue__T_last__T_10_addr] <= buffer_1_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (buffer_1_Queue_reset) begin
      buffer_1_Queue_value <= 1'h0;
    end else if (buffer_1_Queue__T_6) begin
      buffer_1_Queue_value <= buffer_1_Queue__T_12;
    end
    if (buffer_1_Queue_reset) begin
      buffer_1_Queue_value_1 <= 1'h0;
    end else if (buffer_1_Queue__T_8) begin
      buffer_1_Queue_value_1 <= buffer_1_Queue__T_14;
    end
    if (buffer_1_Queue_reset) begin
      buffer_1_Queue__T_1 <= 1'h0;
    end else if (buffer_1_Queue__T_15) begin
      buffer_1_Queue__T_1 <= buffer_1_Queue__T_6;
    end
  end
  always @(posedge buffer_2_Queue_clock) begin
    if(buffer_2_Queue__T_data__T_10_en & buffer_2_Queue__T_data__T_10_mask) begin
      buffer_2_Queue__T_data[buffer_2_Queue__T_data__T_10_addr] <= buffer_2_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(buffer_2_Queue__T_last__T_10_en & buffer_2_Queue__T_last__T_10_mask) begin
      buffer_2_Queue__T_last[buffer_2_Queue__T_last__T_10_addr] <= buffer_2_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (buffer_2_Queue_reset) begin
      buffer_2_Queue_value <= 1'h0;
    end else if (buffer_2_Queue__T_6) begin
      buffer_2_Queue_value <= buffer_2_Queue__T_12;
    end
    if (buffer_2_Queue_reset) begin
      buffer_2_Queue_value_1 <= 1'h0;
    end else if (buffer_2_Queue__T_8) begin
      buffer_2_Queue_value_1 <= buffer_2_Queue__T_14;
    end
    if (buffer_2_Queue_reset) begin
      buffer_2_Queue__T_1 <= 1'h0;
    end else if (buffer_2_Queue__T_15) begin
      buffer_2_Queue__T_1 <= buffer_2_Queue__T_6;
    end
  end
  always @(posedge buffer_3_Queue_clock) begin
    if(buffer_3_Queue__T_data__T_10_en & buffer_3_Queue__T_data__T_10_mask) begin
      buffer_3_Queue__T_data[buffer_3_Queue__T_data__T_10_addr] <= buffer_3_Queue__T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(buffer_3_Queue__T_last__T_10_en & buffer_3_Queue__T_last__T_10_mask) begin
      buffer_3_Queue__T_last[buffer_3_Queue__T_last__T_10_addr] <= buffer_3_Queue__T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (buffer_3_Queue_reset) begin
      buffer_3_Queue_value <= 1'h0;
    end else if (buffer_3_Queue__T_6) begin
      buffer_3_Queue_value <= buffer_3_Queue__T_12;
    end
    if (buffer_3_Queue_reset) begin
      buffer_3_Queue_value_1 <= 1'h0;
    end else if (buffer_3_Queue__T_8) begin
      buffer_3_Queue_value_1 <= buffer_3_Queue__T_14;
    end
    if (buffer_3_Queue_reset) begin
      buffer_3_Queue__T_1 <= 1'h0;
    end else if (buffer_3_Queue__T_15) begin
      buffer_3_Queue__T_1 <= buffer_3_Queue__T_6;
    end
  end
  always @(posedge bus_awIn_0_clock) begin
    if(bus_awIn_0__T__T_10_en & bus_awIn_0__T__T_10_mask) begin
      bus_awIn_0__T[bus_awIn_0__T__T_10_addr] <= bus_awIn_0__T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (bus_awIn_0_reset) begin
      bus_awIn_0_value <= 1'h0;
    end else if (bus_awIn_0__GEN_12) begin
      bus_awIn_0_value <= bus_awIn_0__T_12;
    end
    if (bus_awIn_0_reset) begin
      bus_awIn_0_value_1 <= 1'h0;
    end else if (bus_awIn_0__GEN_11) begin
      bus_awIn_0_value_1 <= bus_awIn_0__T_14;
    end
    if (bus_awIn_0_reset) begin
      bus_awIn_0__T_1 <= 1'h0;
    end else if (bus_awIn_0__T_15) begin
      if (bus_awIn_0__T_4) begin
        if (bus_awIn_0_io_deq_ready) begin
          bus_awIn_0__T_1 <= 1'h0;
        end else begin
          bus_awIn_0__T_1 <= bus_awIn_0__T_6;
        end
      end else begin
        bus_awIn_0__T_1 <= bus_awIn_0__T_6;
      end
    end
  end
  always @(posedge bus_clock) begin
    if (bus_reset) begin
      bus__T_59 <= 3'h0;
    end else begin
      bus__T_59 <= bus__T_64;
    end
    if (bus__T_54) begin
      bus__T_60 <= bus__T_45;
    end
    bus__T_302 <= bus_reset | bus__GEN_18;
    if (bus_reset) begin
      bus__T_373_0 <= 1'h0;
    end else if (bus__T_302) begin
      bus__T_373_0 <= bus__T_344;
    end
    if (bus_reset) begin
      bus__T_373_1 <= 1'h0;
    end else if (bus__T_302) begin
      bus__T_373_1 <= bus__T_345;
    end
    if (bus_reset) begin
      bus__T_373_2 <= 1'h0;
    end else if (bus__T_302) begin
      bus__T_373_2 <= bus__T_346;
    end
    if (bus_reset) begin
      bus__T_313 <= 3'h7;
    end else if (bus__T_330) begin
      bus__T_313 <= bus__T_337;
    end
    if (bus_reset) begin
      bus__T_113 <= 1'h0;
    end else if (bus__T_123) begin
      bus__T_113 <= 1'h0;
    end else begin
      bus__T_113 <= bus__GEN_2;
    end
    if (bus_reset) begin
      bus__T_87 <= 3'h0;
    end else begin
      bus__T_87 <= bus__T_92;
    end
    if (bus__T_83) begin
      bus__T_88 <= bus__T_53;
    end
    bus__T_407 <= bus_reset | bus__GEN_21;
    if (bus_reset) begin
      bus__T_478_0 <= 1'h0;
    end else if (bus__T_407) begin
      bus__T_478_0 <= bus__T_449;
    end
    if (bus_reset) begin
      bus__T_478_1 <= 1'h0;
    end else if (bus__T_407) begin
      bus__T_478_1 <= bus__T_450;
    end
    if (bus_reset) begin
      bus__T_478_2 <= 1'h0;
    end else if (bus__T_407) begin
      bus__T_478_2 <= bus__T_451;
    end
    if (bus_reset) begin
      bus__T_418 <= 3'h7;
    end else if (bus__T_435) begin
      bus__T_418 <= bus__T_442;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_70) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_70) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_76) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_76) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_98) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_98) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_104) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_185) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_185) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_206) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_206) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_229) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_229) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_250) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_250) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_273) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_273) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_294) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_294) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_364) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_364) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_371) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_371) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_469) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_469) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (bus__T_476) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (bus__T_476) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
