module AXI4StreamWidthAdapater_4_to_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [7:0]  auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [7:0] _T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg [1:0] _T_3; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire  _T_4; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire  _T_5; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_6; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_7; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_9; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_10; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_12; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_13; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_15; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_16; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [23:0] _T_18; // @[Cat.scala 29:58]
  wire  ov0; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_20; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_4;
  reg  _T_21; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_5;
  reg  _T_22; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_6;
  reg [1:0] _T_23; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_7;
  wire  _T_25; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_26; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_27; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_29; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_30; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_32; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_33; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_35; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_36; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [3:0] _T_39; // @[Cat.scala 29:58]
  wire  ov1; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_44; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_8;
  wire  _T_46; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_47; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_48; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_8; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov2; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_64; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_9;
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_67; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_68; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_12; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov3; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_84; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_10;
  wire  _T_86; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_87; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_88; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_16; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov4; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  _T_101; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  _T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_104; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_105; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  _T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_108; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_109; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  _T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_112; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_113; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  _T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  _T_116; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_4 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  assign _T_5 = _T_3 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_6 = _T_3 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_7 = _T_5 ? 3'h0 : _T_6; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_0 = _T_4 ? _T_7 : {{1'd0}, _T_3}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_9 = _T_3 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_10 = _T_4 & _T_9; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_12 = _T_3 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_13 = _T_4 & _T_12; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_15 = _T_3 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_16 = _T_4 & _T_15; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_18 = {auto_in_bits_data,_T_2,_T_1}; // @[Cat.scala 29:58]
  assign ov0 = _T_5 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_25 = _T_23 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_26 = _T_23 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_27 = _T_25 ? 3'h0 : _T_26; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_4 = _T_4 ? _T_27 : {{1'd0}, _T_23}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_29 = _T_23 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_30 = _T_4 & _T_29; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_32 = _T_23 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_33 = _T_4 & _T_32; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_35 = _T_23 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_36 = _T_4 & _T_35; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_39 = {auto_in_bits_last,_T_22,_T_21,_T_20}; // @[Cat.scala 29:58]
  assign ov1 = _T_25 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_46 = _T_44 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_47 = _T_44 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_48 = _T_46 ? 3'h0 : _T_47; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_8 = _T_4 ? _T_48 : {{1'd0}, _T_44}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov2 = _T_46 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_66 = _T_64 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_67 = _T_64 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_68 = _T_66 ? 3'h0 : _T_67; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_12 = _T_4 ? _T_68 : {{1'd0}, _T_64}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov3 = _T_66 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_86 = _T_84 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_87 = _T_84 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_88 = _T_86 ? 3'h0 : _T_87; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_16 = _T_4 ? _T_88 : {{1'd0}, _T_84}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov4 = _T_86 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_101 = ov0 == ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  assign _T_103 = _T_101 | reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_104 = ~_T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_105 = ov0 == ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  assign _T_107 = _T_105 | reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_108 = ~_T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_109 = ov0 == ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  assign _T_111 = _T_109 | reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_112 = ~_T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_113 = ov0 == ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  assign _T_115 = _T_113 | reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_116 = ~_T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = _T_5 & auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = {_T_18,_T}; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = _T_39 != 4'h0; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_20 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_22 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_23 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_44 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_64 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_84 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_10) begin
      _T <= auto_in_bits_data;
    end
    if (_T_13) begin
      _T_1 <= auto_in_bits_data;
    end
    if (_T_16) begin
      _T_2 <= auto_in_bits_data;
    end
    if (reset) begin
      _T_3 <= 2'h0;
    end else begin
      _T_3 <= _GEN_0[1:0];
    end
    if (_T_30) begin
      _T_20 <= auto_in_bits_last;
    end
    if (_T_33) begin
      _T_21 <= auto_in_bits_last;
    end
    if (_T_36) begin
      _T_22 <= auto_in_bits_last;
    end
    if (reset) begin
      _T_23 <= 2'h0;
    end else begin
      _T_23 <= _GEN_4[1:0];
    end
    if (reset) begin
      _T_44 <= 2'h0;
    end else begin
      _T_44 <= _GEN_8[1:0];
    end
    if (reset) begin
      _T_64 <= 2'h0;
    end else begin
      _T_64 <= _GEN_12[1:0];
    end
    if (reset) begin
      _T_84 <= 2'h0;
    end else begin
      _T_84 <= _GEN_16[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_104) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_108) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_108) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_112) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_116) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_116) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SDFStageRadix22(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_47; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_49; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_52; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_54; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_56; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_59; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_30; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_32; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_35; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_37; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_39; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_42; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h1; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_47 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_49 = _T_47[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_52 = $signed(_T_49) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_52[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_54 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_56 = _T_54[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_59 = $signed(_T_56) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_59[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_30 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_32 = _T_30[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_35 = $signed(_T_32) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_35[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_37 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_39 = _T_37[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_42 = $signed(_T_39) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_42[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      if (load_input) begin
        feedback_real <= io_in_real;
      end else begin
        feedback_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        feedback_imag <= io_in_imag;
      end else begin
        feedback_imag <= butterfly_outputs_1_imag;
      end
    end
  end
endmodule
module SDFStageRadix22_1(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_50; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_52; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_55; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_57; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_59; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_62; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_33; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_35; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_38; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_40; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_42; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_45; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h2; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_50 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_52 = _T_50[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_55 = $signed(_T_52) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_55[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_57 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_59 = _T_57[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_62 = $signed(_T_59) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_62[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_33 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_35 = _T_33[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_38 = $signed(_T_35) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_38[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_40 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_42 = _T_40[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_45 = $signed(_T_42) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_45[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      feedback_real <= _T_21_real;
    end
    if (io_en) begin
      feedback_imag <= _T_21_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
  end
endmodule
module SDFStageRadix22_2(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_56; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_58; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_61; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_63; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_65; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_68; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_39; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_41; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_44; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_46; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_48; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_51; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h4; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_56 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_58 = _T_56[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_61 = $signed(_T_58) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_61[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_63 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_65 = _T_63[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_68 = $signed(_T_65) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_68[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_39 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_41 = _T_39[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_44 = $signed(_T_41) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_44[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_46 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_48 = _T_46[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_51 = $signed(_T_48) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_51[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      feedback_real <= _T_27_real;
    end
    if (io_en) begin
      feedback_imag <= _T_27_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
  end
endmodule
module SDFStageRadix22_3(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_68; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_70; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_73; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_75; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_77; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_80; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_51; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_53; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_56; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_58; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_60; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_63; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h8; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_68 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_70 = _T_68[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_73 = $signed(_T_70) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_73[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_75 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_77 = _T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_80 = $signed(_T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_80[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_51 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_53 = _T_51[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_56 = $signed(_T_53) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_56[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_58 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_60 = _T_58[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_63 = $signed(_T_60) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_63[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      feedback_real <= _T_39_real;
    end
    if (io_en) begin
      feedback_imag <= _T_39_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
  end
endmodule
module SDFStageRadix22_4(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_92; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_94; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_97; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_99; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_101; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_104; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_75; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_77; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_80; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_82; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_84; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_87; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h10; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_92 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_94 = _T_92[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_97 = $signed(_T_94) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_97[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_99 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_101 = _T_99[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_104 = $signed(_T_101) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_104[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_75 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_77 = _T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_80 = $signed(_T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_80[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_82 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_84 = _T_82[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_87 = $signed(_T_84) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_87[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      feedback_real <= _T_63_real;
    end
    if (io_en) begin
      feedback_imag <= _T_63_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
  end
endmodule
module SDFStageRadix22_5(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_140; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_142; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_145; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_147; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_149; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_152; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [15:0] _T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] _T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] _T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] _T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [15:0] _T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [15:0] _T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [15:0] _T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [15:0] _T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [15:0] _T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [15:0] _T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [15:0] _T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [15:0] _T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [15:0] _T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [15:0] _T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [15:0] _T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [15:0] _T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [15:0] _T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [15:0] _T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [15:0] _T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [15:0] _T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] _T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] _T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] _T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] _T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] _T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [15:0] _T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] _T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] _T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] _T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] _T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_123; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_125; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_128; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_130; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_132; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_135; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h20; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_140 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_142 = _T_140[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_145 = $signed(_T_142) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_145[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_147 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_149 = _T_147[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_152 = $signed(_T_149) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_152[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_123 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_125 = _T_123[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_128 = $signed(_T_125) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_128[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_130 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_132 = _T_130[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_135 = $signed(_T_132) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_135[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_66_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_66_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_69_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_69_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_72_real = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_72_imag = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_75_real = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_75_imag = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_78_real = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_78_imag = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_81_real = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_81_imag = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_84_real = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_84_imag = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_87_real = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_87_imag = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_90_real = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_90_imag = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_93_real = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_93_imag = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_96_real = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_96_imag = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_99_real = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_99_imag = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_102_real = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_102_imag = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_105_real = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_105_imag = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_108_real = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_108_imag = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_111_real = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_111_imag = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      feedback_real <= _T_111_real;
    end
    if (io_en) begin
      feedback_imag <= _T_111_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    if (io_en) begin
      _T_66_real <= _T_63_real;
    end
    if (io_en) begin
      _T_66_imag <= _T_63_imag;
    end
    if (io_en) begin
      _T_69_real <= _T_66_real;
    end
    if (io_en) begin
      _T_69_imag <= _T_66_imag;
    end
    if (io_en) begin
      _T_72_real <= _T_69_real;
    end
    if (io_en) begin
      _T_72_imag <= _T_69_imag;
    end
    if (io_en) begin
      _T_75_real <= _T_72_real;
    end
    if (io_en) begin
      _T_75_imag <= _T_72_imag;
    end
    if (io_en) begin
      _T_78_real <= _T_75_real;
    end
    if (io_en) begin
      _T_78_imag <= _T_75_imag;
    end
    if (io_en) begin
      _T_81_real <= _T_78_real;
    end
    if (io_en) begin
      _T_81_imag <= _T_78_imag;
    end
    if (io_en) begin
      _T_84_real <= _T_81_real;
    end
    if (io_en) begin
      _T_84_imag <= _T_81_imag;
    end
    if (io_en) begin
      _T_87_real <= _T_84_real;
    end
    if (io_en) begin
      _T_87_imag <= _T_84_imag;
    end
    if (io_en) begin
      _T_90_real <= _T_87_real;
    end
    if (io_en) begin
      _T_90_imag <= _T_87_imag;
    end
    if (io_en) begin
      _T_93_real <= _T_90_real;
    end
    if (io_en) begin
      _T_93_imag <= _T_90_imag;
    end
    if (io_en) begin
      _T_96_real <= _T_93_real;
    end
    if (io_en) begin
      _T_96_imag <= _T_93_imag;
    end
    if (io_en) begin
      _T_99_real <= _T_96_real;
    end
    if (io_en) begin
      _T_99_imag <= _T_96_imag;
    end
    if (io_en) begin
      _T_102_real <= _T_99_real;
    end
    if (io_en) begin
      _T_102_imag <= _T_99_imag;
    end
    if (io_en) begin
      _T_105_real <= _T_102_real;
    end
    if (io_en) begin
      _T_105_imag <= _T_102_imag;
    end
    if (io_en) begin
      _T_108_real <= _T_105_real;
    end
    if (io_en) begin
      _T_108_imag <= _T_105_imag;
    end
    if (io_en) begin
      _T_111_real <= _T_108_real;
    end
    if (io_en) begin
      _T_111_imag <= _T_108_imag;
    end
  end
endmodule
module SDFStageRadix22_6(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_236; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_238; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_241; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_243; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_245; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_248; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [15:0] _T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] _T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] _T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] _T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [15:0] _T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [15:0] _T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [15:0] _T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [15:0] _T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [15:0] _T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [15:0] _T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [15:0] _T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [15:0] _T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [15:0] _T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [15:0] _T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [15:0] _T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [15:0] _T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [15:0] _T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [15:0] _T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [15:0] _T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [15:0] _T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] _T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] _T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] _T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] _T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] _T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [15:0] _T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] _T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] _T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] _T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] _T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [15:0] _T_114_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [15:0] _T_114_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [15:0] _T_117_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [15:0] _T_117_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [15:0] _T_120_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [15:0] _T_120_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [15:0] _T_123_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [15:0] _T_123_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [15:0] _T_126_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [15:0] _T_126_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [15:0] _T_129_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [15:0] _T_129_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [15:0] _T_132_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [15:0] _T_132_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [15:0] _T_135_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [15:0] _T_135_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [15:0] _T_138_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [15:0] _T_138_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [15:0] _T_141_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [15:0] _T_141_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [15:0] _T_144_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [15:0] _T_144_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [15:0] _T_147_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [15:0] _T_147_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [15:0] _T_150_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [15:0] _T_150_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [15:0] _T_153_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [15:0] _T_153_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [15:0] _T_156_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [15:0] _T_156_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [15:0] _T_159_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [15:0] _T_159_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [15:0] _T_162_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [15:0] _T_162_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [15:0] _T_165_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [15:0] _T_165_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [15:0] _T_168_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [15:0] _T_168_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [15:0] _T_171_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [15:0] _T_171_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [15:0] _T_174_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [15:0] _T_174_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [15:0] _T_177_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [15:0] _T_177_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [15:0] _T_180_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [15:0] _T_180_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [15:0] _T_183_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [15:0] _T_183_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [15:0] _T_186_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [15:0] _T_186_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [15:0] _T_189_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [15:0] _T_189_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [15:0] _T_192_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [15:0] _T_192_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [15:0] _T_195_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [15:0] _T_195_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [15:0] _T_198_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [15:0] _T_198_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [15:0] _T_201_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [15:0] _T_201_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [15:0] _T_204_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [15:0] _T_204_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [15:0] _T_207_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [15:0] _T_207_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_219; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_221; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_224; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_226; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_228; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_231; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h40; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_236 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_238 = _T_236[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_241 = $signed(_T_238) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_241[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_243 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_245 = _T_243[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_248 = $signed(_T_245) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_248[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_219 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_221 = _T_219[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_224 = $signed(_T_221) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_224[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_226 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_228 = _T_226[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_231 = $signed(_T_228) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_231[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_66_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_66_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_69_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_69_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_72_real = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_72_imag = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_75_real = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_75_imag = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_78_real = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_78_imag = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_81_real = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_81_imag = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_84_real = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_84_imag = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_87_real = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_87_imag = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_90_real = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_90_imag = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_93_real = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_93_imag = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_96_real = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_96_imag = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_99_real = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_99_imag = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_102_real = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_102_imag = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_105_real = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_105_imag = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_108_real = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_108_imag = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_111_real = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_111_imag = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_114_real = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_114_imag = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_117_real = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_117_imag = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_120_real = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_120_imag = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_123_real = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_123_imag = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_126_real = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_126_imag = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_129_real = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_129_imag = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_132_real = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_132_imag = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_135_real = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_135_imag = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_138_real = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_138_imag = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_141_real = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_141_imag = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_144_real = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_144_imag = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_147_real = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_147_imag = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_150_real = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_150_imag = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_153_real = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_153_imag = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_156_real = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_156_imag = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_159_real = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_159_imag = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_162_real = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_162_imag = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_165_real = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_165_imag = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_168_real = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_168_imag = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_171_real = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_171_imag = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_174_real = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_174_imag = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_177_real = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_177_imag = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_180_real = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_180_imag = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_183_real = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_183_imag = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_186_real = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_186_imag = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_189_real = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_189_imag = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_192_real = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_192_imag = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_195_real = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_195_imag = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_198_real = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_198_imag = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_201_real = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_201_imag = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_204_real = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_204_imag = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_207_real = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_207_imag = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      feedback_real <= _T_207_real;
    end
    if (io_en) begin
      feedback_imag <= _T_207_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    if (io_en) begin
      _T_66_real <= _T_63_real;
    end
    if (io_en) begin
      _T_66_imag <= _T_63_imag;
    end
    if (io_en) begin
      _T_69_real <= _T_66_real;
    end
    if (io_en) begin
      _T_69_imag <= _T_66_imag;
    end
    if (io_en) begin
      _T_72_real <= _T_69_real;
    end
    if (io_en) begin
      _T_72_imag <= _T_69_imag;
    end
    if (io_en) begin
      _T_75_real <= _T_72_real;
    end
    if (io_en) begin
      _T_75_imag <= _T_72_imag;
    end
    if (io_en) begin
      _T_78_real <= _T_75_real;
    end
    if (io_en) begin
      _T_78_imag <= _T_75_imag;
    end
    if (io_en) begin
      _T_81_real <= _T_78_real;
    end
    if (io_en) begin
      _T_81_imag <= _T_78_imag;
    end
    if (io_en) begin
      _T_84_real <= _T_81_real;
    end
    if (io_en) begin
      _T_84_imag <= _T_81_imag;
    end
    if (io_en) begin
      _T_87_real <= _T_84_real;
    end
    if (io_en) begin
      _T_87_imag <= _T_84_imag;
    end
    if (io_en) begin
      _T_90_real <= _T_87_real;
    end
    if (io_en) begin
      _T_90_imag <= _T_87_imag;
    end
    if (io_en) begin
      _T_93_real <= _T_90_real;
    end
    if (io_en) begin
      _T_93_imag <= _T_90_imag;
    end
    if (io_en) begin
      _T_96_real <= _T_93_real;
    end
    if (io_en) begin
      _T_96_imag <= _T_93_imag;
    end
    if (io_en) begin
      _T_99_real <= _T_96_real;
    end
    if (io_en) begin
      _T_99_imag <= _T_96_imag;
    end
    if (io_en) begin
      _T_102_real <= _T_99_real;
    end
    if (io_en) begin
      _T_102_imag <= _T_99_imag;
    end
    if (io_en) begin
      _T_105_real <= _T_102_real;
    end
    if (io_en) begin
      _T_105_imag <= _T_102_imag;
    end
    if (io_en) begin
      _T_108_real <= _T_105_real;
    end
    if (io_en) begin
      _T_108_imag <= _T_105_imag;
    end
    if (io_en) begin
      _T_111_real <= _T_108_real;
    end
    if (io_en) begin
      _T_111_imag <= _T_108_imag;
    end
    if (io_en) begin
      _T_114_real <= _T_111_real;
    end
    if (io_en) begin
      _T_114_imag <= _T_111_imag;
    end
    if (io_en) begin
      _T_117_real <= _T_114_real;
    end
    if (io_en) begin
      _T_117_imag <= _T_114_imag;
    end
    if (io_en) begin
      _T_120_real <= _T_117_real;
    end
    if (io_en) begin
      _T_120_imag <= _T_117_imag;
    end
    if (io_en) begin
      _T_123_real <= _T_120_real;
    end
    if (io_en) begin
      _T_123_imag <= _T_120_imag;
    end
    if (io_en) begin
      _T_126_real <= _T_123_real;
    end
    if (io_en) begin
      _T_126_imag <= _T_123_imag;
    end
    if (io_en) begin
      _T_129_real <= _T_126_real;
    end
    if (io_en) begin
      _T_129_imag <= _T_126_imag;
    end
    if (io_en) begin
      _T_132_real <= _T_129_real;
    end
    if (io_en) begin
      _T_132_imag <= _T_129_imag;
    end
    if (io_en) begin
      _T_135_real <= _T_132_real;
    end
    if (io_en) begin
      _T_135_imag <= _T_132_imag;
    end
    if (io_en) begin
      _T_138_real <= _T_135_real;
    end
    if (io_en) begin
      _T_138_imag <= _T_135_imag;
    end
    if (io_en) begin
      _T_141_real <= _T_138_real;
    end
    if (io_en) begin
      _T_141_imag <= _T_138_imag;
    end
    if (io_en) begin
      _T_144_real <= _T_141_real;
    end
    if (io_en) begin
      _T_144_imag <= _T_141_imag;
    end
    if (io_en) begin
      _T_147_real <= _T_144_real;
    end
    if (io_en) begin
      _T_147_imag <= _T_144_imag;
    end
    if (io_en) begin
      _T_150_real <= _T_147_real;
    end
    if (io_en) begin
      _T_150_imag <= _T_147_imag;
    end
    if (io_en) begin
      _T_153_real <= _T_150_real;
    end
    if (io_en) begin
      _T_153_imag <= _T_150_imag;
    end
    if (io_en) begin
      _T_156_real <= _T_153_real;
    end
    if (io_en) begin
      _T_156_imag <= _T_153_imag;
    end
    if (io_en) begin
      _T_159_real <= _T_156_real;
    end
    if (io_en) begin
      _T_159_imag <= _T_156_imag;
    end
    if (io_en) begin
      _T_162_real <= _T_159_real;
    end
    if (io_en) begin
      _T_162_imag <= _T_159_imag;
    end
    if (io_en) begin
      _T_165_real <= _T_162_real;
    end
    if (io_en) begin
      _T_165_imag <= _T_162_imag;
    end
    if (io_en) begin
      _T_168_real <= _T_165_real;
    end
    if (io_en) begin
      _T_168_imag <= _T_165_imag;
    end
    if (io_en) begin
      _T_171_real <= _T_168_real;
    end
    if (io_en) begin
      _T_171_imag <= _T_168_imag;
    end
    if (io_en) begin
      _T_174_real <= _T_171_real;
    end
    if (io_en) begin
      _T_174_imag <= _T_171_imag;
    end
    if (io_en) begin
      _T_177_real <= _T_174_real;
    end
    if (io_en) begin
      _T_177_imag <= _T_174_imag;
    end
    if (io_en) begin
      _T_180_real <= _T_177_real;
    end
    if (io_en) begin
      _T_180_imag <= _T_177_imag;
    end
    if (io_en) begin
      _T_183_real <= _T_180_real;
    end
    if (io_en) begin
      _T_183_imag <= _T_180_imag;
    end
    if (io_en) begin
      _T_186_real <= _T_183_real;
    end
    if (io_en) begin
      _T_186_imag <= _T_183_imag;
    end
    if (io_en) begin
      _T_189_real <= _T_186_real;
    end
    if (io_en) begin
      _T_189_imag <= _T_186_imag;
    end
    if (io_en) begin
      _T_192_real <= _T_189_real;
    end
    if (io_en) begin
      _T_192_imag <= _T_189_imag;
    end
    if (io_en) begin
      _T_195_real <= _T_192_real;
    end
    if (io_en) begin
      _T_195_imag <= _T_192_imag;
    end
    if (io_en) begin
      _T_198_real <= _T_195_real;
    end
    if (io_en) begin
      _T_198_imag <= _T_195_imag;
    end
    if (io_en) begin
      _T_201_real <= _T_198_real;
    end
    if (io_en) begin
      _T_201_imag <= _T_198_imag;
    end
    if (io_en) begin
      _T_204_real <= _T_201_real;
    end
    if (io_en) begin
      _T_204_imag <= _T_201_imag;
    end
    if (io_en) begin
      _T_207_real <= _T_204_real;
    end
    if (io_en) begin
      _T_207_imag <= _T_204_imag;
    end
  end
endmodule
module SDFStageRadix22_7(
  input         clock,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_428; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_430; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_433; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_435; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_437; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_440; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [15:0] _T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] _T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] _T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] _T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [15:0] _T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [15:0] _T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [15:0] _T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [15:0] _T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [15:0] _T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [15:0] _T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [15:0] _T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [15:0] _T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [15:0] _T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [15:0] _T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [15:0] _T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [15:0] _T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [15:0] _T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [15:0] _T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [15:0] _T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [15:0] _T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] _T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] _T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] _T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] _T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] _T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [15:0] _T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] _T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] _T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] _T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] _T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [15:0] _T_114_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [15:0] _T_114_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [15:0] _T_117_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [15:0] _T_117_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [15:0] _T_120_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [15:0] _T_120_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [15:0] _T_123_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [15:0] _T_123_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [15:0] _T_126_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [15:0] _T_126_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [15:0] _T_129_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [15:0] _T_129_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [15:0] _T_132_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [15:0] _T_132_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [15:0] _T_135_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [15:0] _T_135_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [15:0] _T_138_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [15:0] _T_138_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [15:0] _T_141_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [15:0] _T_141_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [15:0] _T_144_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [15:0] _T_144_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [15:0] _T_147_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [15:0] _T_147_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [15:0] _T_150_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [15:0] _T_150_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [15:0] _T_153_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [15:0] _T_153_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [15:0] _T_156_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [15:0] _T_156_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [15:0] _T_159_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [15:0] _T_159_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [15:0] _T_162_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [15:0] _T_162_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [15:0] _T_165_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [15:0] _T_165_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [15:0] _T_168_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [15:0] _T_168_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [15:0] _T_171_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [15:0] _T_171_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [15:0] _T_174_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [15:0] _T_174_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [15:0] _T_177_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [15:0] _T_177_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [15:0] _T_180_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [15:0] _T_180_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [15:0] _T_183_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [15:0] _T_183_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [15:0] _T_186_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [15:0] _T_186_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [15:0] _T_189_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [15:0] _T_189_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [15:0] _T_192_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [15:0] _T_192_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [15:0] _T_195_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [15:0] _T_195_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [15:0] _T_198_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [15:0] _T_198_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [15:0] _T_201_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [15:0] _T_201_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [15:0] _T_204_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [15:0] _T_204_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [15:0] _T_207_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [15:0] _T_207_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [15:0] _T_210_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [15:0] _T_210_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [15:0] _T_213_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [15:0] _T_213_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [15:0] _T_216_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [15:0] _T_216_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [15:0] _T_219_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [15:0] _T_219_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [15:0] _T_222_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [15:0] _T_222_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [15:0] _T_225_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [15:0] _T_225_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [15:0] _T_228_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [15:0] _T_228_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [15:0] _T_231_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [15:0] _T_231_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [15:0] _T_234_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [15:0] _T_234_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [15:0] _T_237_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [15:0] _T_237_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [15:0] _T_240_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [15:0] _T_240_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [15:0] _T_243_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [15:0] _T_243_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [15:0] _T_246_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [15:0] _T_246_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [15:0] _T_249_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [15:0] _T_249_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [15:0] _T_252_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [15:0] _T_252_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [15:0] _T_255_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [15:0] _T_255_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [15:0] _T_258_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [15:0] _T_258_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [15:0] _T_261_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [15:0] _T_261_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [15:0] _T_264_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [15:0] _T_264_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [15:0] _T_267_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [15:0] _T_267_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [15:0] _T_270_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [15:0] _T_270_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [15:0] _T_273_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [15:0] _T_273_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [15:0] _T_276_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [15:0] _T_276_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [15:0] _T_279_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [15:0] _T_279_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [15:0] _T_282_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [15:0] _T_282_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [15:0] _T_285_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [15:0] _T_285_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [15:0] _T_288_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [15:0] _T_288_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [15:0] _T_291_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [15:0] _T_291_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [15:0] _T_294_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [15:0] _T_294_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [15:0] _T_297_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [15:0] _T_297_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [15:0] _T_300_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [15:0] _T_300_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [15:0] _T_303_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [15:0] _T_303_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [15:0] _T_306_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [15:0] _T_306_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [15:0] _T_309_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [15:0] _T_309_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [15:0] _T_312_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [15:0] _T_312_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [15:0] _T_315_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [15:0] _T_315_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [15:0] _T_318_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [15:0] _T_318_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [15:0] _T_321_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [15:0] _T_321_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [15:0] _T_324_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [15:0] _T_324_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [15:0] _T_327_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [15:0] _T_327_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [15:0] _T_330_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [15:0] _T_330_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [15:0] _T_333_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [15:0] _T_333_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [15:0] _T_336_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [15:0] _T_336_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [15:0] _T_339_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [15:0] _T_339_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [15:0] _T_342_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [15:0] _T_342_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [15:0] _T_345_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [15:0] _T_345_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [15:0] _T_348_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [15:0] _T_348_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [15:0] _T_351_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [15:0] _T_351_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [15:0] _T_354_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [15:0] _T_354_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [15:0] _T_357_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [15:0] _T_357_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [15:0] _T_360_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [15:0] _T_360_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [15:0] _T_363_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [15:0] _T_363_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [15:0] _T_366_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [15:0] _T_366_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [15:0] _T_369_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [15:0] _T_369_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [15:0] _T_372_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [15:0] _T_372_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [15:0] _T_375_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [15:0] _T_375_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [15:0] _T_378_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [15:0] _T_378_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [15:0] _T_381_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [15:0] _T_381_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [15:0] _T_384_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [15:0] _T_384_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [15:0] _T_387_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [15:0] _T_387_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [15:0] _T_390_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [15:0] _T_390_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [15:0] _T_393_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [15:0] _T_393_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [15:0] _T_396_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [15:0] _T_396_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [15:0] _T_399_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [15:0] _T_399_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_411; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_413; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_416; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_418; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_420; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_423; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  assign load_input = io_cntr < 9'h80; // @[UIntTypeClass.scala 52:47]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_428 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_430 = _T_428[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_433 = $signed(_T_430) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_433[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_435 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_437 = _T_435[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_440 = $signed(_T_437) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_440[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_411 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_413 = _T_411[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_416 = $signed(_T_413) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_416[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_418 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_420 = _T_418[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_423 = $signed(_T_420) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_423[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  feedback_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  feedback_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_66_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_66_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_69_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_69_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_72_real = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_72_imag = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_75_real = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_75_imag = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_78_real = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_78_imag = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_81_real = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_81_imag = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_84_real = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_84_imag = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_87_real = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_87_imag = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_90_real = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_90_imag = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_93_real = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_93_imag = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_96_real = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_96_imag = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_99_real = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_99_imag = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_102_real = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_102_imag = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_105_real = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_105_imag = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_108_real = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_108_imag = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_111_real = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_111_imag = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_114_real = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_114_imag = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_117_real = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_117_imag = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_120_real = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_120_imag = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_123_real = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_123_imag = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_126_real = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_126_imag = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_129_real = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_129_imag = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_132_real = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_132_imag = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_135_real = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_135_imag = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_138_real = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_138_imag = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_141_real = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_141_imag = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_144_real = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_144_imag = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_147_real = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_147_imag = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_150_real = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_150_imag = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_153_real = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_153_imag = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_156_real = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_156_imag = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_159_real = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_159_imag = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_162_real = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_162_imag = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_165_real = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_165_imag = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_168_real = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_168_imag = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_171_real = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_171_imag = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_174_real = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_174_imag = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_177_real = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_177_imag = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_180_real = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_180_imag = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_183_real = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_183_imag = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_186_real = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_186_imag = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_189_real = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_189_imag = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_192_real = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_192_imag = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_195_real = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_195_imag = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_198_real = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_198_imag = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_201_real = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_201_imag = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_204_real = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_204_imag = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_207_real = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_207_imag = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_210_real = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_210_imag = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_213_real = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_213_imag = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_216_real = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_216_imag = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_219_real = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_219_imag = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_222_real = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_222_imag = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_225_real = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_225_imag = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_228_real = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_228_imag = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_231_real = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_231_imag = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_234_real = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_234_imag = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_237_real = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_237_imag = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_240_real = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_240_imag = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_243_real = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_243_imag = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_246_real = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_246_imag = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_249_real = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_249_imag = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_252_real = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_252_imag = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_255_real = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_255_imag = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_258_real = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_258_imag = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_261_real = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_261_imag = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_264_real = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_264_imag = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_267_real = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_267_imag = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_270_real = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_270_imag = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_273_real = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_273_imag = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_276_real = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_276_imag = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_279_real = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_279_imag = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_282_real = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_282_imag = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_285_real = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_285_imag = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_288_real = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_288_imag = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_291_real = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_291_imag = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_294_real = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_294_imag = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_297_real = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_297_imag = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_300_real = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_300_imag = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_303_real = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_303_imag = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_306_real = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_306_imag = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_309_real = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_309_imag = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_312_real = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_312_imag = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_315_real = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_315_imag = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_318_real = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_318_imag = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_321_real = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_321_imag = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_324_real = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_324_imag = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_327_real = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_327_imag = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_330_real = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_330_imag = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_333_real = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_333_imag = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_336_real = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_336_imag = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_339_real = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_339_imag = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_342_real = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_342_imag = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_345_real = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_345_imag = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_348_real = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_348_imag = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_351_real = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_351_imag = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_354_real = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_354_imag = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_357_real = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_357_imag = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_360_real = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_360_imag = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_363_real = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_363_imag = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_366_real = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_366_imag = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_369_real = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_369_imag = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_372_real = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_372_imag = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_375_real = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_375_imag = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_378_real = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_378_imag = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_381_real = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_381_imag = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_384_real = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_384_imag = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_387_real = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_387_imag = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_390_real = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_390_imag = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_393_real = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_393_imag = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_396_real = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_396_imag = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_399_real = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_399_imag = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      feedback_real <= _T_399_real;
    end
    if (io_en) begin
      feedback_imag <= _T_399_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    if (io_en) begin
      _T_66_real <= _T_63_real;
    end
    if (io_en) begin
      _T_66_imag <= _T_63_imag;
    end
    if (io_en) begin
      _T_69_real <= _T_66_real;
    end
    if (io_en) begin
      _T_69_imag <= _T_66_imag;
    end
    if (io_en) begin
      _T_72_real <= _T_69_real;
    end
    if (io_en) begin
      _T_72_imag <= _T_69_imag;
    end
    if (io_en) begin
      _T_75_real <= _T_72_real;
    end
    if (io_en) begin
      _T_75_imag <= _T_72_imag;
    end
    if (io_en) begin
      _T_78_real <= _T_75_real;
    end
    if (io_en) begin
      _T_78_imag <= _T_75_imag;
    end
    if (io_en) begin
      _T_81_real <= _T_78_real;
    end
    if (io_en) begin
      _T_81_imag <= _T_78_imag;
    end
    if (io_en) begin
      _T_84_real <= _T_81_real;
    end
    if (io_en) begin
      _T_84_imag <= _T_81_imag;
    end
    if (io_en) begin
      _T_87_real <= _T_84_real;
    end
    if (io_en) begin
      _T_87_imag <= _T_84_imag;
    end
    if (io_en) begin
      _T_90_real <= _T_87_real;
    end
    if (io_en) begin
      _T_90_imag <= _T_87_imag;
    end
    if (io_en) begin
      _T_93_real <= _T_90_real;
    end
    if (io_en) begin
      _T_93_imag <= _T_90_imag;
    end
    if (io_en) begin
      _T_96_real <= _T_93_real;
    end
    if (io_en) begin
      _T_96_imag <= _T_93_imag;
    end
    if (io_en) begin
      _T_99_real <= _T_96_real;
    end
    if (io_en) begin
      _T_99_imag <= _T_96_imag;
    end
    if (io_en) begin
      _T_102_real <= _T_99_real;
    end
    if (io_en) begin
      _T_102_imag <= _T_99_imag;
    end
    if (io_en) begin
      _T_105_real <= _T_102_real;
    end
    if (io_en) begin
      _T_105_imag <= _T_102_imag;
    end
    if (io_en) begin
      _T_108_real <= _T_105_real;
    end
    if (io_en) begin
      _T_108_imag <= _T_105_imag;
    end
    if (io_en) begin
      _T_111_real <= _T_108_real;
    end
    if (io_en) begin
      _T_111_imag <= _T_108_imag;
    end
    if (io_en) begin
      _T_114_real <= _T_111_real;
    end
    if (io_en) begin
      _T_114_imag <= _T_111_imag;
    end
    if (io_en) begin
      _T_117_real <= _T_114_real;
    end
    if (io_en) begin
      _T_117_imag <= _T_114_imag;
    end
    if (io_en) begin
      _T_120_real <= _T_117_real;
    end
    if (io_en) begin
      _T_120_imag <= _T_117_imag;
    end
    if (io_en) begin
      _T_123_real <= _T_120_real;
    end
    if (io_en) begin
      _T_123_imag <= _T_120_imag;
    end
    if (io_en) begin
      _T_126_real <= _T_123_real;
    end
    if (io_en) begin
      _T_126_imag <= _T_123_imag;
    end
    if (io_en) begin
      _T_129_real <= _T_126_real;
    end
    if (io_en) begin
      _T_129_imag <= _T_126_imag;
    end
    if (io_en) begin
      _T_132_real <= _T_129_real;
    end
    if (io_en) begin
      _T_132_imag <= _T_129_imag;
    end
    if (io_en) begin
      _T_135_real <= _T_132_real;
    end
    if (io_en) begin
      _T_135_imag <= _T_132_imag;
    end
    if (io_en) begin
      _T_138_real <= _T_135_real;
    end
    if (io_en) begin
      _T_138_imag <= _T_135_imag;
    end
    if (io_en) begin
      _T_141_real <= _T_138_real;
    end
    if (io_en) begin
      _T_141_imag <= _T_138_imag;
    end
    if (io_en) begin
      _T_144_real <= _T_141_real;
    end
    if (io_en) begin
      _T_144_imag <= _T_141_imag;
    end
    if (io_en) begin
      _T_147_real <= _T_144_real;
    end
    if (io_en) begin
      _T_147_imag <= _T_144_imag;
    end
    if (io_en) begin
      _T_150_real <= _T_147_real;
    end
    if (io_en) begin
      _T_150_imag <= _T_147_imag;
    end
    if (io_en) begin
      _T_153_real <= _T_150_real;
    end
    if (io_en) begin
      _T_153_imag <= _T_150_imag;
    end
    if (io_en) begin
      _T_156_real <= _T_153_real;
    end
    if (io_en) begin
      _T_156_imag <= _T_153_imag;
    end
    if (io_en) begin
      _T_159_real <= _T_156_real;
    end
    if (io_en) begin
      _T_159_imag <= _T_156_imag;
    end
    if (io_en) begin
      _T_162_real <= _T_159_real;
    end
    if (io_en) begin
      _T_162_imag <= _T_159_imag;
    end
    if (io_en) begin
      _T_165_real <= _T_162_real;
    end
    if (io_en) begin
      _T_165_imag <= _T_162_imag;
    end
    if (io_en) begin
      _T_168_real <= _T_165_real;
    end
    if (io_en) begin
      _T_168_imag <= _T_165_imag;
    end
    if (io_en) begin
      _T_171_real <= _T_168_real;
    end
    if (io_en) begin
      _T_171_imag <= _T_168_imag;
    end
    if (io_en) begin
      _T_174_real <= _T_171_real;
    end
    if (io_en) begin
      _T_174_imag <= _T_171_imag;
    end
    if (io_en) begin
      _T_177_real <= _T_174_real;
    end
    if (io_en) begin
      _T_177_imag <= _T_174_imag;
    end
    if (io_en) begin
      _T_180_real <= _T_177_real;
    end
    if (io_en) begin
      _T_180_imag <= _T_177_imag;
    end
    if (io_en) begin
      _T_183_real <= _T_180_real;
    end
    if (io_en) begin
      _T_183_imag <= _T_180_imag;
    end
    if (io_en) begin
      _T_186_real <= _T_183_real;
    end
    if (io_en) begin
      _T_186_imag <= _T_183_imag;
    end
    if (io_en) begin
      _T_189_real <= _T_186_real;
    end
    if (io_en) begin
      _T_189_imag <= _T_186_imag;
    end
    if (io_en) begin
      _T_192_real <= _T_189_real;
    end
    if (io_en) begin
      _T_192_imag <= _T_189_imag;
    end
    if (io_en) begin
      _T_195_real <= _T_192_real;
    end
    if (io_en) begin
      _T_195_imag <= _T_192_imag;
    end
    if (io_en) begin
      _T_198_real <= _T_195_real;
    end
    if (io_en) begin
      _T_198_imag <= _T_195_imag;
    end
    if (io_en) begin
      _T_201_real <= _T_198_real;
    end
    if (io_en) begin
      _T_201_imag <= _T_198_imag;
    end
    if (io_en) begin
      _T_204_real <= _T_201_real;
    end
    if (io_en) begin
      _T_204_imag <= _T_201_imag;
    end
    if (io_en) begin
      _T_207_real <= _T_204_real;
    end
    if (io_en) begin
      _T_207_imag <= _T_204_imag;
    end
    if (io_en) begin
      _T_210_real <= _T_207_real;
    end
    if (io_en) begin
      _T_210_imag <= _T_207_imag;
    end
    if (io_en) begin
      _T_213_real <= _T_210_real;
    end
    if (io_en) begin
      _T_213_imag <= _T_210_imag;
    end
    if (io_en) begin
      _T_216_real <= _T_213_real;
    end
    if (io_en) begin
      _T_216_imag <= _T_213_imag;
    end
    if (io_en) begin
      _T_219_real <= _T_216_real;
    end
    if (io_en) begin
      _T_219_imag <= _T_216_imag;
    end
    if (io_en) begin
      _T_222_real <= _T_219_real;
    end
    if (io_en) begin
      _T_222_imag <= _T_219_imag;
    end
    if (io_en) begin
      _T_225_real <= _T_222_real;
    end
    if (io_en) begin
      _T_225_imag <= _T_222_imag;
    end
    if (io_en) begin
      _T_228_real <= _T_225_real;
    end
    if (io_en) begin
      _T_228_imag <= _T_225_imag;
    end
    if (io_en) begin
      _T_231_real <= _T_228_real;
    end
    if (io_en) begin
      _T_231_imag <= _T_228_imag;
    end
    if (io_en) begin
      _T_234_real <= _T_231_real;
    end
    if (io_en) begin
      _T_234_imag <= _T_231_imag;
    end
    if (io_en) begin
      _T_237_real <= _T_234_real;
    end
    if (io_en) begin
      _T_237_imag <= _T_234_imag;
    end
    if (io_en) begin
      _T_240_real <= _T_237_real;
    end
    if (io_en) begin
      _T_240_imag <= _T_237_imag;
    end
    if (io_en) begin
      _T_243_real <= _T_240_real;
    end
    if (io_en) begin
      _T_243_imag <= _T_240_imag;
    end
    if (io_en) begin
      _T_246_real <= _T_243_real;
    end
    if (io_en) begin
      _T_246_imag <= _T_243_imag;
    end
    if (io_en) begin
      _T_249_real <= _T_246_real;
    end
    if (io_en) begin
      _T_249_imag <= _T_246_imag;
    end
    if (io_en) begin
      _T_252_real <= _T_249_real;
    end
    if (io_en) begin
      _T_252_imag <= _T_249_imag;
    end
    if (io_en) begin
      _T_255_real <= _T_252_real;
    end
    if (io_en) begin
      _T_255_imag <= _T_252_imag;
    end
    if (io_en) begin
      _T_258_real <= _T_255_real;
    end
    if (io_en) begin
      _T_258_imag <= _T_255_imag;
    end
    if (io_en) begin
      _T_261_real <= _T_258_real;
    end
    if (io_en) begin
      _T_261_imag <= _T_258_imag;
    end
    if (io_en) begin
      _T_264_real <= _T_261_real;
    end
    if (io_en) begin
      _T_264_imag <= _T_261_imag;
    end
    if (io_en) begin
      _T_267_real <= _T_264_real;
    end
    if (io_en) begin
      _T_267_imag <= _T_264_imag;
    end
    if (io_en) begin
      _T_270_real <= _T_267_real;
    end
    if (io_en) begin
      _T_270_imag <= _T_267_imag;
    end
    if (io_en) begin
      _T_273_real <= _T_270_real;
    end
    if (io_en) begin
      _T_273_imag <= _T_270_imag;
    end
    if (io_en) begin
      _T_276_real <= _T_273_real;
    end
    if (io_en) begin
      _T_276_imag <= _T_273_imag;
    end
    if (io_en) begin
      _T_279_real <= _T_276_real;
    end
    if (io_en) begin
      _T_279_imag <= _T_276_imag;
    end
    if (io_en) begin
      _T_282_real <= _T_279_real;
    end
    if (io_en) begin
      _T_282_imag <= _T_279_imag;
    end
    if (io_en) begin
      _T_285_real <= _T_282_real;
    end
    if (io_en) begin
      _T_285_imag <= _T_282_imag;
    end
    if (io_en) begin
      _T_288_real <= _T_285_real;
    end
    if (io_en) begin
      _T_288_imag <= _T_285_imag;
    end
    if (io_en) begin
      _T_291_real <= _T_288_real;
    end
    if (io_en) begin
      _T_291_imag <= _T_288_imag;
    end
    if (io_en) begin
      _T_294_real <= _T_291_real;
    end
    if (io_en) begin
      _T_294_imag <= _T_291_imag;
    end
    if (io_en) begin
      _T_297_real <= _T_294_real;
    end
    if (io_en) begin
      _T_297_imag <= _T_294_imag;
    end
    if (io_en) begin
      _T_300_real <= _T_297_real;
    end
    if (io_en) begin
      _T_300_imag <= _T_297_imag;
    end
    if (io_en) begin
      _T_303_real <= _T_300_real;
    end
    if (io_en) begin
      _T_303_imag <= _T_300_imag;
    end
    if (io_en) begin
      _T_306_real <= _T_303_real;
    end
    if (io_en) begin
      _T_306_imag <= _T_303_imag;
    end
    if (io_en) begin
      _T_309_real <= _T_306_real;
    end
    if (io_en) begin
      _T_309_imag <= _T_306_imag;
    end
    if (io_en) begin
      _T_312_real <= _T_309_real;
    end
    if (io_en) begin
      _T_312_imag <= _T_309_imag;
    end
    if (io_en) begin
      _T_315_real <= _T_312_real;
    end
    if (io_en) begin
      _T_315_imag <= _T_312_imag;
    end
    if (io_en) begin
      _T_318_real <= _T_315_real;
    end
    if (io_en) begin
      _T_318_imag <= _T_315_imag;
    end
    if (io_en) begin
      _T_321_real <= _T_318_real;
    end
    if (io_en) begin
      _T_321_imag <= _T_318_imag;
    end
    if (io_en) begin
      _T_324_real <= _T_321_real;
    end
    if (io_en) begin
      _T_324_imag <= _T_321_imag;
    end
    if (io_en) begin
      _T_327_real <= _T_324_real;
    end
    if (io_en) begin
      _T_327_imag <= _T_324_imag;
    end
    if (io_en) begin
      _T_330_real <= _T_327_real;
    end
    if (io_en) begin
      _T_330_imag <= _T_327_imag;
    end
    if (io_en) begin
      _T_333_real <= _T_330_real;
    end
    if (io_en) begin
      _T_333_imag <= _T_330_imag;
    end
    if (io_en) begin
      _T_336_real <= _T_333_real;
    end
    if (io_en) begin
      _T_336_imag <= _T_333_imag;
    end
    if (io_en) begin
      _T_339_real <= _T_336_real;
    end
    if (io_en) begin
      _T_339_imag <= _T_336_imag;
    end
    if (io_en) begin
      _T_342_real <= _T_339_real;
    end
    if (io_en) begin
      _T_342_imag <= _T_339_imag;
    end
    if (io_en) begin
      _T_345_real <= _T_342_real;
    end
    if (io_en) begin
      _T_345_imag <= _T_342_imag;
    end
    if (io_en) begin
      _T_348_real <= _T_345_real;
    end
    if (io_en) begin
      _T_348_imag <= _T_345_imag;
    end
    if (io_en) begin
      _T_351_real <= _T_348_real;
    end
    if (io_en) begin
      _T_351_imag <= _T_348_imag;
    end
    if (io_en) begin
      _T_354_real <= _T_351_real;
    end
    if (io_en) begin
      _T_354_imag <= _T_351_imag;
    end
    if (io_en) begin
      _T_357_real <= _T_354_real;
    end
    if (io_en) begin
      _T_357_imag <= _T_354_imag;
    end
    if (io_en) begin
      _T_360_real <= _T_357_real;
    end
    if (io_en) begin
      _T_360_imag <= _T_357_imag;
    end
    if (io_en) begin
      _T_363_real <= _T_360_real;
    end
    if (io_en) begin
      _T_363_imag <= _T_360_imag;
    end
    if (io_en) begin
      _T_366_real <= _T_363_real;
    end
    if (io_en) begin
      _T_366_imag <= _T_363_imag;
    end
    if (io_en) begin
      _T_369_real <= _T_366_real;
    end
    if (io_en) begin
      _T_369_imag <= _T_366_imag;
    end
    if (io_en) begin
      _T_372_real <= _T_369_real;
    end
    if (io_en) begin
      _T_372_imag <= _T_369_imag;
    end
    if (io_en) begin
      _T_375_real <= _T_372_real;
    end
    if (io_en) begin
      _T_375_imag <= _T_372_imag;
    end
    if (io_en) begin
      _T_378_real <= _T_375_real;
    end
    if (io_en) begin
      _T_378_imag <= _T_375_imag;
    end
    if (io_en) begin
      _T_381_real <= _T_378_real;
    end
    if (io_en) begin
      _T_381_imag <= _T_378_imag;
    end
    if (io_en) begin
      _T_384_real <= _T_381_real;
    end
    if (io_en) begin
      _T_384_imag <= _T_381_imag;
    end
    if (io_en) begin
      _T_387_real <= _T_384_real;
    end
    if (io_en) begin
      _T_387_imag <= _T_384_imag;
    end
    if (io_en) begin
      _T_390_real <= _T_387_real;
    end
    if (io_en) begin
      _T_390_imag <= _T_387_imag;
    end
    if (io_en) begin
      _T_393_real <= _T_390_real;
    end
    if (io_en) begin
      _T_393_imag <= _T_390_imag;
    end
    if (io_en) begin
      _T_396_real <= _T_393_real;
    end
    if (io_en) begin
      _T_396_imag <= _T_393_imag;
    end
    if (io_en) begin
      _T_399_real <= _T_396_real;
    end
    if (io_en) begin
      _T_399_imag <= _T_396_imag;
    end
  end
endmodule
module SDFStageRadix22_8(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [8:0]  io_cntr,
  input         io_en
);
  wire [7:0] SRAM_depth_256_width_32_mem_R0_addr; // @[ShiftRegisterMem.scala 48:28]
  wire  SRAM_depth_256_width_32_mem_R0_en; // @[ShiftRegisterMem.scala 48:28]
  wire  SRAM_depth_256_width_32_mem_R0_clk; // @[ShiftRegisterMem.scala 48:28]
  wire [15:0] SRAM_depth_256_width_32_mem_R0_data_real; // @[ShiftRegisterMem.scala 48:28]
  wire [15:0] SRAM_depth_256_width_32_mem_R0_data_imag; // @[ShiftRegisterMem.scala 48:28]
  wire [7:0] SRAM_depth_256_width_32_mem_W0_addr; // @[ShiftRegisterMem.scala 48:28]
  wire  SRAM_depth_256_width_32_mem_W0_en; // @[ShiftRegisterMem.scala 48:28]
  wire  SRAM_depth_256_width_32_mem_W0_clk; // @[ShiftRegisterMem.scala 48:28]
  wire [15:0] SRAM_depth_256_width_32_mem_W0_data_real; // @[ShiftRegisterMem.scala 48:28]
  wire [15:0] SRAM_depth_256_width_32_mem_W0_data_imag; // @[ShiftRegisterMem.scala 48:28]
  wire  load_input; // @[UIntTypeClass.scala 52:47]
  wire [15:0] feedback_real; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_57; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_59; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_62; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  wire [15:0] feedback_imag; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_64; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_66; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_69; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [7:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [7:0] _T_22; // @[Counter.scala 39:22]
  reg [7:0] _T_26; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_40; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_42; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_45; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_real; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _T_47; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_49; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_52; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butt_out_0_imag; // @[FixedPointTypeClass.scala 176:41]
  SRAM_depth_256_width_32_mem SRAM_depth_256_width_32_mem ( // @[ShiftRegisterMem.scala 48:28]
    .R0_addr(SRAM_depth_256_width_32_mem_R0_addr),
    .R0_en(SRAM_depth_256_width_32_mem_R0_en),
    .R0_clk(SRAM_depth_256_width_32_mem_R0_clk),
    .R0_data_real(SRAM_depth_256_width_32_mem_R0_data_real),
    .R0_data_imag(SRAM_depth_256_width_32_mem_R0_data_imag),
    .W0_addr(SRAM_depth_256_width_32_mem_W0_addr),
    .W0_en(SRAM_depth_256_width_32_mem_W0_en),
    .W0_clk(SRAM_depth_256_width_32_mem_W0_clk),
    .W0_data_real(SRAM_depth_256_width_32_mem_W0_data_real),
    .W0_data_imag(SRAM_depth_256_width_32_mem_W0_data_imag)
  );
  assign load_input = io_cntr < 9'h100; // @[UIntTypeClass.scala 52:47]
  assign feedback_real = SRAM_depth_256_width_32_mem_R0_data_real; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  assign butt_outputs_1_real = $signed(feedback_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_57 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_59 = _T_57[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_62 = $signed(_T_59) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_62[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign feedback_imag = SRAM_depth_256_width_32_mem_R0_data_imag; // @[SDFChainRadix22.scala 470:23 SDFChainRadix22.scala 483:17]
  assign butt_outputs_1_imag = $signed(feedback_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_64 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_66 = _T_64[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_69 = $signed(_T_66) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_69[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_22 = value + 8'h1; // @[Counter.scala 39:22]
  assign butt_outputs_0_real = $signed(feedback_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(feedback_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_40 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_42 = _T_40[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_45 = $signed(_T_42) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_real = _T_45[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_47 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_49 = _T_47[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_52 = $signed(_T_49) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butt_out_0_imag = _T_52[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign io_out_real = load_input ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 463:10]
  assign io_out_imag = load_input ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 463:10]
  assign SRAM_depth_256_width_32_mem_R0_addr = value; // @[ShiftRegisterMem.scala 53:25]
  assign SRAM_depth_256_width_32_mem_R0_en = io_en; // @[ShiftRegisterMem.scala 48:28 Counter.scala 39:13]
  assign SRAM_depth_256_width_32_mem_R0_clk = clock; // @[ShiftRegisterMem.scala 53:25]
  assign SRAM_depth_256_width_32_mem_W0_addr = _T_26;
  assign SRAM_depth_256_width_32_mem_W0_en = io_en; // @[ShiftRegisterMem.scala 48:28]
  assign SRAM_depth_256_width_32_mem_W0_clk = clock;
  assign SRAM_depth_256_width_32_mem_W0_data_real = load_input ? $signed(io_in_real) : $signed(butterfly_outputs_1_real);
  assign SRAM_depth_256_width_32_mem_W0_data_imag = load_input ? $signed(io_in_imag) : $signed(butterfly_outputs_1_imag);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 8'h0;
    end else if (io_en) begin
      value <= _T_22;
    end
    if (reset) begin
      _T_26 <= 8'hff;
    end else if (io_en) begin
      _T_26 <= value;
    end
  end
endmodule
module SDFChainRadix22(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  output        io_lastOut,
  input         io_lastIn,
  output        io_busy
);
  wire  sdf_stages_0_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_0_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_0_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_0_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_0_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_0_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_0_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_1_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_1_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_1_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_1_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_1_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_1_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_1_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_2_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_2_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_2_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_2_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_2_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_2_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_2_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_3_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_3_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_3_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_3_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_3_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_3_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_3_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_4_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_4_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_4_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_4_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_4_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_4_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_4_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_5_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_5_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_5_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_5_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_5_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_5_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_5_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_6_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_6_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_6_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_6_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_6_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_6_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_6_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_7_clock; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_7_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_7_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_7_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_7_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_7_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_7_io_en; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_8_clock; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_8_reset; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_8_io_in_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_8_io_in_imag; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_8_io_out_real; // @[SDFChainRadix22.scala 164:25]
  wire [15:0] sdf_stages_8_io_out_imag; // @[SDFChainRadix22.scala 164:25]
  wire [8:0] sdf_stages_8_io_cntr; // @[SDFChainRadix22.scala 164:25]
  wire  sdf_stages_8_io_en; // @[SDFChainRadix22.scala 164:25]
  reg [1:0] state; // @[SDFChainRadix22.scala 56:22]
  reg [31:0] _RAND_0;
  reg  initialOutDone; // @[SDFChainRadix22.scala 59:31]
  reg [31:0] _RAND_1;
  reg [9:0] cnt; // @[SDFChainRadix22.scala 60:20]
  reg [31:0] _RAND_2;
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  fireLast; // @[SDFChainRadix22.scala 79:28]
  wire [8:0] _T_48; // @[SDFChainRadix22.scala 81:45]
  wire  _T_53; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_0; // @[SDFChainRadix22.scala 90:27]
  wire  _T_56; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1; // @[SDFChainRadix22.scala 93:23]
  wire  _T_57; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_2; // @[SDFChainRadix22.scala 98:25]
  wire [1:0] _GEN_3; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67]
  wire [1:0] state_next; // @[Conditional.scala 40:58]
  reg [8:0] cntValidOut; // @[SDFChainRadix22.scala 106:28]
  reg [31:0] _RAND_3;
  wire [9:0] _T_59; // @[SDFChainRadix22.scala 111:44]
  wire [9:0] _GEN_2109; // @[SDFChainRadix22.scala 111:29]
  wire  _T_60; // @[SDFChainRadix22.scala 111:29]
  wire  _T_61; // @[Decoupled.scala 40:37]
  wire  pktEnd; // @[SDFChainRadix22.scala 111:52]
  wire  _T_62; // @[SDFChainRadix22.scala 114:20]
  wire [8:0] cntr_wires_0; // @[SDFChainRadix22.scala 52:24 SDFChainRadix22.scala 185:29]
  wire [8:0] _GEN_20; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] _GEN_21; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] _GEN_22; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] _GEN_23; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] _GEN_24; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] _GEN_25; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] _GEN_26; // @[SDFChainRadix22.scala 126:79]
  wire [8:0] _GEN_27; // @[SDFChainRadix22.scala 126:79]
  wire [9:0] _GEN_2110; // @[SDFChainRadix22.scala 126:79]
  wire  _T_76; // @[SDFChainRadix22.scala 130:31]
  wire  _T_77; // @[SDFChainRadix22.scala 130:42]
  wire [8:0] _T_80; // @[SDFChainRadix22.scala 134:32]
  wire  _T_83; // @[SDFChainRadix22.scala 144:90]
  wire  _T_122; // @[SDFChainRadix22.scala 173:54]
  wire  enableInit; // @[SDFChainRadix22.scala 173:33]
  wire [9:0] _T_125; // @[SDFChainRadix22.scala 179:16]
  wire [9:0] _T_145; // @[SDFChainRadix22.scala 193:37]
  wire  _T_146; // @[SDFChainRadix22.scala 193:22]
  wire  _T_147; // @[SDFChainRadix22.scala 193:44]
  wire  _GEN_45; // @[SDFChainRadix22.scala 196:36]
  wire  _GEN_46; // @[SDFChainRadix22.scala 193:60]
  wire [8:0] _T_166; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_171; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] _T_173; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_178; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] _T_180; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_185; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] _T_187; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_192; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] _T_194; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_199; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] _T_201; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_206; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] _T_208; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_213; // @[SDFChainRadix22.scala 224:68]
  wire [8:0] _T_215; // @[SDFChainRadix22.scala 224:38]
  wire [8:0] _T_220; // @[SDFChainRadix22.scala 224:68]
  wire [1:0] _GEN_52; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] _GEN_53; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] _GEN_54; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] _GEN_55; // @[SDFChainRadix22.scala 291:27]
  wire [1:0] _GEN_56; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_59; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_60; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_61; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_62; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_63; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] twiddles_1_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] _T_261; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] outputWires_0_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  wire [15:0] outputWires_0_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  wire [16:0] _T_262; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] _T_263; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] _GEN_2112; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_264; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2113; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_265; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2114; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_266; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] _T_267; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] _T_268; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] _T_274; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_275; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] _T_278; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_279; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_286; // @[SDFChainRadix22.scala 328:32]
  wire  _T_287; // @[SDFChainRadix22.scala 328:78]
  wire  _T_288; // @[SDFChainRadix22.scala 328:65]
  wire  _T_289; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] outputWires_1_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] _T_295; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] outputWires_1_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [3:0] _GEN_82; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_83; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_84; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_85; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_86; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_87; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_88; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_89; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_90; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_91; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_92; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_93; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_94; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_95; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_96; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_97; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_98; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_99; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_100; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_101; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_102; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_103; // @[SDFChainRadix22.scala 291:27]
  wire [3:0] _GEN_104; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_107; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_108; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_109; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_110; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_111; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_112; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_113; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_114; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_115; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_116; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_117; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_118; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_119; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_120; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_121; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_122; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_123; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_124; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_125; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_126; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_127; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_128; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_129; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_130; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_131; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_132; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_133; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_134; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_135; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] twiddles_3_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] _T_393; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] outputWires_2_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] outputWires_2_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [16:0] _T_394; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] _T_395; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] _GEN_2115; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_396; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2116; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_397; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2117; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_398; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] _T_399; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] _T_400; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] _T_406; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_407; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] _T_410; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_411; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_418; // @[SDFChainRadix22.scala 328:32]
  wire  _T_419; // @[SDFChainRadix22.scala 328:78]
  wire  _T_420; // @[SDFChainRadix22.scala 328:65]
  wire  _T_421; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] outputWires_3_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] _T_427; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] outputWires_3_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [5:0] _GEN_202; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_203; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_204; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_205; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_206; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_207; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_208; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_209; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_210; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_211; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_212; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_213; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_214; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_215; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_216; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_217; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_218; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_219; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_220; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_221; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_222; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_223; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_224; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_225; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_226; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_227; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_228; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_229; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_230; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_231; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_232; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_233; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_234; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_235; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_236; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_237; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_238; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_239; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_240; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_241; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_242; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_243; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_244; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_245; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_246; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_247; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_248; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_249; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_250; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_251; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_252; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_253; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_254; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_255; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_256; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_257; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_258; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_259; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_260; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_261; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_262; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_263; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_264; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_265; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_266; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_267; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_268; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_269; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_270; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_271; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_272; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_273; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_274; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_275; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_276; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_277; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_278; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_279; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_280; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_281; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_282; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_283; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_284; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_285; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_286; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_287; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_288; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_289; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_290; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_291; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_292; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_293; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_294; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_295; // @[SDFChainRadix22.scala 291:27]
  wire [5:0] _GEN_296; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_299; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_300; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_301; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_302; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_303; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_304; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_305; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_306; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_307; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_308; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_309; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_310; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_311; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_312; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_313; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_314; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_315; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_316; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_317; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_318; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_319; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_320; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_321; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_322; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_323; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_324; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_325; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_326; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_327; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_328; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_329; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_330; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_331; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_332; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_333; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_334; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_335; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_336; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_337; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_338; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_339; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_340; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_341; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_342; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_343; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_344; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_345; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_346; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_347; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_348; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_349; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_350; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_351; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_352; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_353; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_354; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_355; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_356; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_357; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_358; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_359; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_360; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_361; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_362; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_363; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_364; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_365; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_366; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_367; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_368; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_369; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_370; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_371; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_372; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_373; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_374; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_375; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_376; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_377; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_378; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_379; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_380; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_381; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_382; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_383; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_384; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_385; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_386; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_387; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_388; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_389; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_390; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_391; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_392; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_393; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_394; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_395; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_396; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_397; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_398; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_399; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_400; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_401; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_402; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_403; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_404; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_405; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_406; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_407; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_408; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_409; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_410; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_411; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_412; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_413; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_414; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_415; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_416; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_417; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_418; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_419; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_420; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_421; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_422; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_423; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] twiddles_5_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] _T_765; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] outputWires_4_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] outputWires_4_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [16:0] _T_766; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] _T_767; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] _GEN_2118; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_768; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2119; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_769; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2120; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_770; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] _T_771; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] _T_772; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] _T_778; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_779; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] _T_782; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_783; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_790; // @[SDFChainRadix22.scala 328:32]
  wire  _T_791; // @[SDFChainRadix22.scala 328:78]
  wire  _T_792; // @[SDFChainRadix22.scala 328:65]
  wire  _T_793; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] outputWires_5_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] _T_799; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] outputWires_5_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [7:0] _GEN_682; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_683; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_684; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_685; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_686; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_687; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_688; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_689; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_690; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_691; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_692; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_693; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_694; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_695; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_696; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_697; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_698; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_699; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_700; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_701; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_702; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_703; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_704; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_705; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_706; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_707; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_708; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_709; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_710; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_711; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_712; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_713; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_714; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_715; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_716; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_717; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_718; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_719; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_720; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_721; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_722; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_723; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_724; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_725; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_726; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_727; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_728; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_729; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_730; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_731; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_732; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_733; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_734; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_735; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_736; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_737; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_738; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_739; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_740; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_741; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_742; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_743; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_744; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_745; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_746; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_747; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_748; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_749; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_750; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_751; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_752; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_753; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_754; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_755; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_756; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_757; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_758; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_759; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_760; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_761; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_762; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_763; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_764; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_765; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_766; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_767; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_768; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_769; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_770; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_771; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_772; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_773; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_774; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_775; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_776; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_777; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_778; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_779; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_780; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_781; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_782; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_783; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_784; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_785; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_786; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_787; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_788; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_789; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_790; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_791; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_792; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_793; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_794; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_795; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_796; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_797; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_798; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_799; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_800; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_801; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_802; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_803; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_804; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_805; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_806; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_807; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_808; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_809; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_810; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_811; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_812; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_813; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_814; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_815; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_816; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_817; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_818; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_819; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_820; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_821; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_822; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_823; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_824; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_825; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_826; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_827; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_828; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_829; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_830; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_831; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_832; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_833; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_834; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_835; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_836; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_837; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_838; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_839; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_840; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_841; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_842; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_843; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_844; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_845; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_846; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_847; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_848; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_849; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_850; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_851; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_852; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_853; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_854; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_855; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_856; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_857; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_858; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_859; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_860; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_861; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_862; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_863; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_864; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_865; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_866; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_867; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_868; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_869; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_870; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_871; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_872; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_873; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_874; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_875; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_876; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_877; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_878; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_879; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_880; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_881; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_882; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_883; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_884; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_885; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_886; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_887; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_888; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_889; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_890; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_891; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_892; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_893; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_894; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_895; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_896; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_897; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_898; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_899; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_900; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_901; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_902; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_903; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_904; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_905; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_906; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_907; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_908; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_909; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_910; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_911; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_912; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_913; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_914; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_915; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_916; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_917; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_918; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_919; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_920; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_921; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_922; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_923; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_924; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_925; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_926; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_927; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_928; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_929; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_930; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_931; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_932; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_933; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_934; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_935; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_936; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_937; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_938; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_939; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_940; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_941; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_942; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_943; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_944; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_945; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_946; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_947; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_948; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_949; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_950; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_951; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_952; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_953; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_954; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_955; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_956; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_957; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_958; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_959; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_960; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_961; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_962; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_963; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_964; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_965; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_966; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_967; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_968; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_969; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_970; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_971; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_972; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_973; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_974; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_975; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_976; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_977; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_978; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_979; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_980; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_981; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_982; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_983; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_984; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_985; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_986; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_987; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_988; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_989; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_990; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_991; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_992; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_993; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_994; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_995; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_996; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_997; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_998; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_999; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1000; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1001; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1002; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1003; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1004; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1005; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1006; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1007; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1008; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1009; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1010; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1011; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1012; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1013; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1014; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1015; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1016; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1017; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1018; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1019; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1020; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1021; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1022; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1023; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1024; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1025; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1026; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1027; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1028; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1029; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1030; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1031; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1032; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1033; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1034; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1035; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1036; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1037; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1038; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1039; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1040; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1041; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1042; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1043; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1044; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1045; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1046; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1047; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1048; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1049; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1050; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1051; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1052; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1053; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1054; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1055; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1056; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1057; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1058; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1059; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1060; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1061; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1062; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1063; // @[SDFChainRadix22.scala 291:27]
  wire [7:0] _GEN_1064; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1067; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1068; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1069; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1070; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1071; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1072; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1073; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1074; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1075; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1076; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1077; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1078; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1079; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1080; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1081; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1082; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1083; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1084; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1085; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1086; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1087; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1088; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1089; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1090; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1091; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1092; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1093; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1094; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1095; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1096; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1097; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1098; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1099; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1100; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1101; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1102; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1103; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1104; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1105; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1106; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1107; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1108; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1109; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1110; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1111; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1112; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1113; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1114; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1115; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1116; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1117; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1118; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1119; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1120; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1121; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1122; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1123; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1124; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1125; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1126; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1127; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1128; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1129; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1130; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1131; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1132; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1133; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1134; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1135; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1136; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1137; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1138; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1139; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1140; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1141; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1142; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1143; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1144; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1145; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1146; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1147; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1148; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1149; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1150; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1151; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1152; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1153; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1154; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1155; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1156; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1157; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1158; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1159; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1160; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1161; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1162; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1163; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1164; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1165; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1166; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1167; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1168; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1169; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1170; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1171; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1172; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1173; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1174; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1175; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1176; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1177; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1178; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1179; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1180; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1181; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1182; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1183; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1184; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1185; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1186; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1187; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1188; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1189; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1190; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1191; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1192; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1193; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1194; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1195; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1196; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1197; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1198; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1199; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1200; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1201; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1202; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1203; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1204; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1205; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1206; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1207; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1208; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1209; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1210; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1211; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1212; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1213; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1214; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1215; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1216; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1217; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1218; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1219; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1220; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1221; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1222; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1223; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1224; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1225; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1226; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1227; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1228; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1229; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1230; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1231; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1232; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1233; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1234; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1235; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1236; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1237; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1238; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1239; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1240; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1241; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1242; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1243; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1244; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1245; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1246; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1247; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1248; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1249; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1250; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1251; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1252; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1253; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1254; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1255; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1256; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1257; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1258; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1259; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1260; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1261; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1262; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1263; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1264; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1265; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1266; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1267; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1268; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1269; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1270; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1271; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1272; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1273; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1274; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1275; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1276; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1277; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1278; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1279; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1280; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1281; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1282; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1283; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1284; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1285; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1286; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1287; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1288; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1289; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1290; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1291; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1292; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1293; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1294; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1295; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1296; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1297; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1298; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1299; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1300; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1301; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1302; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1303; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1304; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1305; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1306; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1307; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1308; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1309; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1310; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1311; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1312; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1313; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1314; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1315; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1316; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1317; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1318; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1319; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1320; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1321; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1322; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1323; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1324; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1325; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1326; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1327; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1328; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1329; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1330; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1331; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1332; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1333; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1334; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1335; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1336; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1337; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1338; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1339; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1340; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1341; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1342; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1343; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1344; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1345; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1346; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1347; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1348; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1349; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1350; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1351; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1352; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1353; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1354; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1355; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1356; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1357; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1358; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1359; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1360; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1361; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1362; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1363; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1364; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1365; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1366; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1367; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1368; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1369; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1370; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1371; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1372; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1373; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1374; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1375; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1376; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1377; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1378; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1379; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1380; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1381; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1382; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1383; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1384; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1385; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1386; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1387; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1388; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1389; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1390; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1391; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1392; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1393; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1394; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1395; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1396; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1397; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1398; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1399; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1400; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1401; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1402; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1403; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1404; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1405; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1406; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1407; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1408; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1409; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1410; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1411; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1412; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1413; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1414; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1415; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1416; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1417; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1418; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1419; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1420; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1421; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1422; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1423; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1424; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1425; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1426; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1427; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1428; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1429; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1430; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1431; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1432; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1433; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1434; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1435; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1436; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1437; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1438; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1439; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1440; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1441; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1442; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1443; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1444; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1445; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1446; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1447; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1448; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1449; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1450; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1451; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1452; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1453; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1454; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1455; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1456; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1457; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1458; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1459; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1460; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1461; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1462; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1463; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1464; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1465; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1466; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1467; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1468; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1469; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1470; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1471; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1472; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1473; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1474; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1475; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1476; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1477; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1478; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1479; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1480; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1481; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1482; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1483; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1484; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1485; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1486; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1487; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1488; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1489; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1490; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1491; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1492; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1493; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1494; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1495; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1496; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1497; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1498; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1499; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1500; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1501; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1502; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1503; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1504; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1505; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1506; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1507; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1508; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1509; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1510; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1511; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1512; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1513; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1514; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1515; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1516; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1517; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1518; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1519; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1520; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1521; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1522; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1523; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1524; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1525; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1526; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1527; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1528; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1529; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1530; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1531; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1532; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1533; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1534; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1535; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1536; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1537; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1538; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1539; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1540; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1541; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1542; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1543; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1544; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1545; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1546; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1547; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1548; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1549; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1550; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1551; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1552; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1553; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1554; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1555; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1556; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1557; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1558; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1559; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1560; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1561; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1562; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1563; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1564; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1565; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1566; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1567; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1568; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1569; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1570; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1571; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1572; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1573; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1574; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] _GEN_1575; // @[SDFChainRadix22.scala 291:27]
  wire [15:0] twiddles_7_imag; // @[SDFChainRadix22.scala 291:27]
  wire [16:0] _T_2096; // @[FixedPointTypeClass.scala 24:22]
  wire [15:0] outputWires_6_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] outputWires_6_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [16:0] _T_2097; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] _T_2098; // @[FixedPointTypeClass.scala 33:22]
  wire [16:0] _GEN_2121; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_2099; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2122; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_2100; // @[FixedPointTypeClass.scala 211:35]
  wire [16:0] _GEN_2123; // @[FixedPointTypeClass.scala 211:35]
  wire [32:0] _T_2101; // @[FixedPointTypeClass.scala 211:35]
  wire [33:0] _T_2102; // @[FixedPointTypeClass.scala 33:22]
  wire [33:0] _T_2103; // @[FixedPointTypeClass.scala 24:22]
  wire [33:0] _T_2109; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_2110; // @[FixedPointTypeClass.scala 176:41]
  wire [33:0] _T_2113; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_2114; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_2121; // @[SDFChainRadix22.scala 328:32]
  wire  _T_2122; // @[SDFChainRadix22.scala 328:78]
  wire  _T_2123; // @[SDFChainRadix22.scala 328:65]
  wire  _T_2124; // @[SDFChainRadix22.scala 328:19]
  wire [15:0] outputWires_7_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] _T_2130; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] outputWires_7_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  wire [15:0] _GEN_2091; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2092; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2093; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2094; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2095; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2096; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2097; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2098; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2099; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2100; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2101; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2102; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2103; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] _GEN_2104; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] outputWires_8_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] _GEN_2105; // @[SDFChainRadix22.scala 364:24]
  wire [15:0] outputWires_8_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  wire [15:0] _GEN_2106; // @[SDFChainRadix22.scala 364:24]
  wire  _T_2140; // @[SDFChainRadix22.scala 368:33]
  wire  _T_2141; // @[SDFChainRadix22.scala 368:127]
  wire  _T_2142; // @[SDFChainRadix22.scala 368:117]
  wire [29:0] _GEN_2124; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] _GEN_2107; // @[SDFChainRadix22.scala 375:33]
  wire [29:0] _GEN_2125; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] _GEN_2108; // @[SDFChainRadix22.scala 375:33]
  wire [17:0] _GEN_2126; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 396:27]
  wire [17:0] _GEN_2128; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 397:27]
  SDFStageRadix22 sdf_stages_0 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_0_clock),
    .io_in_real(sdf_stages_0_io_in_real),
    .io_in_imag(sdf_stages_0_io_in_imag),
    .io_out_real(sdf_stages_0_io_out_real),
    .io_out_imag(sdf_stages_0_io_out_imag),
    .io_cntr(sdf_stages_0_io_cntr),
    .io_en(sdf_stages_0_io_en)
  );
  SDFStageRadix22_1 sdf_stages_1 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_1_clock),
    .io_in_real(sdf_stages_1_io_in_real),
    .io_in_imag(sdf_stages_1_io_in_imag),
    .io_out_real(sdf_stages_1_io_out_real),
    .io_out_imag(sdf_stages_1_io_out_imag),
    .io_cntr(sdf_stages_1_io_cntr),
    .io_en(sdf_stages_1_io_en)
  );
  SDFStageRadix22_2 sdf_stages_2 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_2_clock),
    .io_in_real(sdf_stages_2_io_in_real),
    .io_in_imag(sdf_stages_2_io_in_imag),
    .io_out_real(sdf_stages_2_io_out_real),
    .io_out_imag(sdf_stages_2_io_out_imag),
    .io_cntr(sdf_stages_2_io_cntr),
    .io_en(sdf_stages_2_io_en)
  );
  SDFStageRadix22_3 sdf_stages_3 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_3_clock),
    .io_in_real(sdf_stages_3_io_in_real),
    .io_in_imag(sdf_stages_3_io_in_imag),
    .io_out_real(sdf_stages_3_io_out_real),
    .io_out_imag(sdf_stages_3_io_out_imag),
    .io_cntr(sdf_stages_3_io_cntr),
    .io_en(sdf_stages_3_io_en)
  );
  SDFStageRadix22_4 sdf_stages_4 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_4_clock),
    .io_in_real(sdf_stages_4_io_in_real),
    .io_in_imag(sdf_stages_4_io_in_imag),
    .io_out_real(sdf_stages_4_io_out_real),
    .io_out_imag(sdf_stages_4_io_out_imag),
    .io_cntr(sdf_stages_4_io_cntr),
    .io_en(sdf_stages_4_io_en)
  );
  SDFStageRadix22_5 sdf_stages_5 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_5_clock),
    .io_in_real(sdf_stages_5_io_in_real),
    .io_in_imag(sdf_stages_5_io_in_imag),
    .io_out_real(sdf_stages_5_io_out_real),
    .io_out_imag(sdf_stages_5_io_out_imag),
    .io_cntr(sdf_stages_5_io_cntr),
    .io_en(sdf_stages_5_io_en)
  );
  SDFStageRadix22_6 sdf_stages_6 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_6_clock),
    .io_in_real(sdf_stages_6_io_in_real),
    .io_in_imag(sdf_stages_6_io_in_imag),
    .io_out_real(sdf_stages_6_io_out_real),
    .io_out_imag(sdf_stages_6_io_out_imag),
    .io_cntr(sdf_stages_6_io_cntr),
    .io_en(sdf_stages_6_io_en)
  );
  SDFStageRadix22_7 sdf_stages_7 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_7_clock),
    .io_in_real(sdf_stages_7_io_in_real),
    .io_in_imag(sdf_stages_7_io_in_imag),
    .io_out_real(sdf_stages_7_io_out_real),
    .io_out_imag(sdf_stages_7_io_out_imag),
    .io_cntr(sdf_stages_7_io_cntr),
    .io_en(sdf_stages_7_io_en)
  );
  SDFStageRadix22_8 sdf_stages_8 ( // @[SDFChainRadix22.scala 164:25]
    .clock(sdf_stages_8_clock),
    .reset(sdf_stages_8_reset),
    .io_in_real(sdf_stages_8_io_in_real),
    .io_in_imag(sdf_stages_8_io_in_imag),
    .io_out_real(sdf_stages_8_io_out_real),
    .io_out_imag(sdf_stages_8_io_out_imag),
    .io_cntr(sdf_stages_8_io_cntr),
    .io_en(sdf_stages_8_io_en)
  );
  assign _T_46 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign fireLast = io_lastIn & _T_46; // @[SDFChainRadix22.scala 79:28]
  assign _T_48 = 9'h9 - 9'h1; // @[SDFChainRadix22.scala 81:45]
  assign _T_53 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_0 = _T_46 ? 2'h1 : state; // @[SDFChainRadix22.scala 90:27]
  assign _T_56 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _GEN_1 = fireLast ? 2'h2 : state; // @[SDFChainRadix22.scala 93:23]
  assign _T_57 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_2 = io_lastOut ? 2'h0 : state; // @[SDFChainRadix22.scala 98:25]
  assign _GEN_3 = _T_57 ? _GEN_2 : state; // @[Conditional.scala 39:67]
  assign _GEN_4 = _T_56 ? _GEN_1 : _GEN_3; // @[Conditional.scala 39:67]
  assign state_next = _T_53 ? _GEN_0 : _GEN_4; // @[Conditional.scala 40:58]
  assign _T_59 = 10'h200 - 10'h1; // @[SDFChainRadix22.scala 111:44]
  assign _GEN_2109 = {{1'd0}, cntValidOut}; // @[SDFChainRadix22.scala 111:29]
  assign _T_60 = _GEN_2109 == _T_59; // @[SDFChainRadix22.scala 111:29]
  assign _T_61 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign pktEnd = _T_60 & _T_61; // @[SDFChainRadix22.scala 111:52]
  assign _T_62 = state_next == 2'h0; // @[SDFChainRadix22.scala 114:20]
  assign cntr_wires_0 = cnt[8:0]; // @[SDFChainRadix22.scala 52:24 SDFChainRadix22.scala 185:29]
  assign _GEN_20 = 4'h1 == _T_48[3:0] ? cntr_wires_0 : cntr_wires_0; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_21 = 4'h2 == _T_48[3:0] ? cntr_wires_0 : _GEN_20; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_22 = 4'h3 == _T_48[3:0] ? cntr_wires_0 : _GEN_21; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_23 = 4'h4 == _T_48[3:0] ? cntr_wires_0 : _GEN_22; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_24 = 4'h5 == _T_48[3:0] ? cntr_wires_0 : _GEN_23; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_25 = 4'h6 == _T_48[3:0] ? cntr_wires_0 : _GEN_24; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_26 = 4'h7 == _T_48[3:0] ? cntr_wires_0 : _GEN_25; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_27 = 4'h8 == _T_48[3:0] ? cntr_wires_0 : _GEN_26; // @[SDFChainRadix22.scala 126:79]
  assign _GEN_2110 = {{1'd0}, _GEN_27}; // @[SDFChainRadix22.scala 126:79]
  assign _T_76 = _T_62 & pktEnd; // @[SDFChainRadix22.scala 130:31]
  assign _T_77 = _T_76 | pktEnd; // @[SDFChainRadix22.scala 130:42]
  assign _T_80 = cntValidOut + 9'h1; // @[SDFChainRadix22.scala 134:32]
  assign _T_83 = state == 2'h2; // @[SDFChainRadix22.scala 144:90]
  assign _T_122 = _T_83 & io_out_ready; // @[SDFChainRadix22.scala 173:54]
  assign enableInit = _T_46 | _T_122; // @[SDFChainRadix22.scala 173:33]
  assign _T_125 = cnt + 10'h1; // @[SDFChainRadix22.scala 179:16]
  assign _T_145 = 10'h200 - 10'h2; // @[SDFChainRadix22.scala 193:37]
  assign _T_146 = _GEN_2110 == _T_145; // @[SDFChainRadix22.scala 193:22]
  assign _T_147 = _T_146 & enableInit; // @[SDFChainRadix22.scala 193:44]
  assign _GEN_45 = _T_62 ? 1'h0 : initialOutDone; // @[SDFChainRadix22.scala 196:36]
  assign _GEN_46 = _T_147 | _GEN_45; // @[SDFChainRadix22.scala 193:60]
  assign _T_166 = cntr_wires_0 - 9'h0; // @[SDFChainRadix22.scala 224:38]
  assign _T_171 = 9'h1 - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _T_173 = cntr_wires_0 - _T_171; // @[SDFChainRadix22.scala 224:38]
  assign _T_178 = 9'h3 - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _T_180 = cntr_wires_0 - _T_178; // @[SDFChainRadix22.scala 224:38]
  assign _T_185 = 9'h7 - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _T_187 = cntr_wires_0 - _T_185; // @[SDFChainRadix22.scala 224:38]
  assign _T_192 = 9'hf - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _T_194 = cntr_wires_0 - _T_192; // @[SDFChainRadix22.scala 224:38]
  assign _T_199 = 9'h1f - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _T_201 = cntr_wires_0 - _T_199; // @[SDFChainRadix22.scala 224:38]
  assign _T_206 = 9'h3f - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _T_208 = cntr_wires_0 - _T_206; // @[SDFChainRadix22.scala 224:38]
  assign _T_213 = 9'h7f - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _T_215 = cntr_wires_0 - _T_213; // @[SDFChainRadix22.scala 224:38]
  assign _T_220 = 9'hff - 9'h0; // @[SDFChainRadix22.scala 224:68]
  assign _GEN_52 = 3'h3 == _T_173[2:0] ? 2'h2 : 2'h0; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_53 = 3'h4 == _T_173[2:0] ? 2'h0 : _GEN_52; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_54 = 3'h5 == _T_173[2:0] ? 2'h1 : _GEN_53; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_55 = 3'h6 == _T_173[2:0] ? 2'h0 : _GEN_54; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_56 = 3'h7 == _T_173[2:0] ? 2'h3 : _GEN_55; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_59 = 2'h1 == _GEN_56 ? $signed(16'sh2d41) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_60 = 2'h1 == _GEN_56 ? $signed(-16'sh2d41) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_61 = 2'h2 == _GEN_56 ? $signed(16'sh0) : $signed(_GEN_59); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_62 = 2'h2 == _GEN_56 ? $signed(-16'sh4000) : $signed(_GEN_60); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_63 = 2'h3 == _GEN_56 ? $signed(-16'sh2d41) : $signed(_GEN_61); // @[SDFChainRadix22.scala 291:27]
  assign twiddles_1_imag = 2'h3 == _GEN_56 ? $signed(-16'sh2d41) : $signed(_GEN_62); // @[SDFChainRadix22.scala 291:27]
  assign _T_261 = $signed(_GEN_63) + $signed(twiddles_1_imag); // @[FixedPointTypeClass.scala 24:22]
  assign outputWires_0_real = sdf_stages_0_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  assign outputWires_0_imag = sdf_stages_0_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 348:32]
  assign _T_262 = $signed(outputWires_0_real) + $signed(outputWires_0_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_263 = $signed(outputWires_0_imag) - $signed(outputWires_0_real); // @[FixedPointTypeClass.scala 33:22]
  assign _GEN_2112 = {{1{outputWires_0_real[15]}},outputWires_0_real}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_264 = $signed(_GEN_2112) * $signed(_T_261); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2113 = {{1{twiddles_1_imag[15]}},twiddles_1_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_265 = $signed(_T_262) * $signed(_GEN_2113); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2114 = {{1{_GEN_63[15]}},_GEN_63}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_266 = $signed(_T_263) * $signed(_GEN_2114); // @[FixedPointTypeClass.scala 211:35]
  assign _T_267 = $signed(_T_264) - $signed(_T_265); // @[FixedPointTypeClass.scala 33:22]
  assign _T_268 = $signed(_T_264) + $signed(_T_266); // @[FixedPointTypeClass.scala 24:22]
  assign _T_274 = $signed(_T_267) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_275 = _T_274[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_278 = $signed(_T_268) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_279 = _T_278[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_286 = sdf_stages_2_io_cntr < 9'h4; // @[SDFChainRadix22.scala 328:32]
  assign _T_287 = sdf_stages_2_io_cntr < 9'h6; // @[SDFChainRadix22.scala 328:78]
  assign _T_288 = _T_287 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign _T_289 = _T_286 ? 1'h0 : _T_288; // @[SDFChainRadix22.scala 328:19]
  assign outputWires_1_real = sdf_stages_1_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _T_295 = 16'sh0 - $signed(outputWires_1_real); // @[FixedPointTypeClass.scala 39:43]
  assign outputWires_1_imag = sdf_stages_1_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _GEN_82 = 5'h9 == _T_187[4:0] ? 4'h2 : 4'h0; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_83 = 5'ha == _T_187[4:0] ? 4'h4 : _GEN_82; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_84 = 5'hb == _T_187[4:0] ? 4'h6 : _GEN_83; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_85 = 5'hc == _T_187[4:0] ? 4'h8 : _GEN_84; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_86 = 5'hd == _T_187[4:0] ? 4'ha : _GEN_85; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_87 = 5'he == _T_187[4:0] ? 4'hb : _GEN_86; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_88 = 5'hf == _T_187[4:0] ? 4'hc : _GEN_87; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_89 = 5'h10 == _T_187[4:0] ? 4'h0 : _GEN_88; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_90 = 5'h11 == _T_187[4:0] ? 4'h1 : _GEN_89; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_91 = 5'h12 == _T_187[4:0] ? 4'h2 : _GEN_90; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_92 = 5'h13 == _T_187[4:0] ? 4'h3 : _GEN_91; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_93 = 5'h14 == _T_187[4:0] ? 4'h4 : _GEN_92; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_94 = 5'h15 == _T_187[4:0] ? 4'h5 : _GEN_93; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_95 = 5'h16 == _T_187[4:0] ? 4'h6 : _GEN_94; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_96 = 5'h17 == _T_187[4:0] ? 4'h7 : _GEN_95; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_97 = 5'h18 == _T_187[4:0] ? 4'h0 : _GEN_96; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_98 = 5'h19 == _T_187[4:0] ? 4'h3 : _GEN_97; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_99 = 5'h1a == _T_187[4:0] ? 4'h6 : _GEN_98; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_100 = 5'h1b == _T_187[4:0] ? 4'h9 : _GEN_99; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_101 = 5'h1c == _T_187[4:0] ? 4'hb : _GEN_100; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_102 = 5'h1d == _T_187[4:0] ? 4'hd : _GEN_101; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_103 = 5'h1e == _T_187[4:0] ? 4'he : _GEN_102; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_104 = 5'h1f == _T_187[4:0] ? 4'hf : _GEN_103; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_107 = 4'h1 == _GEN_104 ? $signed(16'sh3ec5) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_108 = 4'h1 == _GEN_104 ? $signed(-16'shc7c) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_109 = 4'h2 == _GEN_104 ? $signed(16'sh3b21) : $signed(_GEN_107); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_110 = 4'h2 == _GEN_104 ? $signed(-16'sh187e) : $signed(_GEN_108); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_111 = 4'h3 == _GEN_104 ? $signed(16'sh3537) : $signed(_GEN_109); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_112 = 4'h3 == _GEN_104 ? $signed(-16'sh238e) : $signed(_GEN_110); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_113 = 4'h4 == _GEN_104 ? $signed(16'sh2d41) : $signed(_GEN_111); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_114 = 4'h4 == _GEN_104 ? $signed(-16'sh2d41) : $signed(_GEN_112); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_115 = 4'h5 == _GEN_104 ? $signed(16'sh238e) : $signed(_GEN_113); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_116 = 4'h5 == _GEN_104 ? $signed(-16'sh3537) : $signed(_GEN_114); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_117 = 4'h6 == _GEN_104 ? $signed(16'sh187e) : $signed(_GEN_115); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_118 = 4'h6 == _GEN_104 ? $signed(-16'sh3b21) : $signed(_GEN_116); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_119 = 4'h7 == _GEN_104 ? $signed(16'shc7c) : $signed(_GEN_117); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_120 = 4'h7 == _GEN_104 ? $signed(-16'sh3ec5) : $signed(_GEN_118); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_121 = 4'h8 == _GEN_104 ? $signed(16'sh0) : $signed(_GEN_119); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_122 = 4'h8 == _GEN_104 ? $signed(-16'sh4000) : $signed(_GEN_120); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_123 = 4'h9 == _GEN_104 ? $signed(-16'shc7c) : $signed(_GEN_121); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_124 = 4'h9 == _GEN_104 ? $signed(-16'sh3ec5) : $signed(_GEN_122); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_125 = 4'ha == _GEN_104 ? $signed(-16'sh187e) : $signed(_GEN_123); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_126 = 4'ha == _GEN_104 ? $signed(-16'sh3b21) : $signed(_GEN_124); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_127 = 4'hb == _GEN_104 ? $signed(-16'sh2d41) : $signed(_GEN_125); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_128 = 4'hb == _GEN_104 ? $signed(-16'sh2d41) : $signed(_GEN_126); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_129 = 4'hc == _GEN_104 ? $signed(-16'sh3b21) : $signed(_GEN_127); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_130 = 4'hc == _GEN_104 ? $signed(-16'sh187e) : $signed(_GEN_128); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_131 = 4'hd == _GEN_104 ? $signed(-16'sh3ec5) : $signed(_GEN_129); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_132 = 4'hd == _GEN_104 ? $signed(-16'shc7c) : $signed(_GEN_130); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_133 = 4'he == _GEN_104 ? $signed(-16'sh3b21) : $signed(_GEN_131); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_134 = 4'he == _GEN_104 ? $signed(16'sh187e) : $signed(_GEN_132); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_135 = 4'hf == _GEN_104 ? $signed(-16'sh238e) : $signed(_GEN_133); // @[SDFChainRadix22.scala 291:27]
  assign twiddles_3_imag = 4'hf == _GEN_104 ? $signed(16'sh3537) : $signed(_GEN_134); // @[SDFChainRadix22.scala 291:27]
  assign _T_393 = $signed(_GEN_135) + $signed(twiddles_3_imag); // @[FixedPointTypeClass.scala 24:22]
  assign outputWires_2_real = sdf_stages_2_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign outputWires_2_imag = sdf_stages_2_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign _T_394 = $signed(outputWires_2_real) + $signed(outputWires_2_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_395 = $signed(outputWires_2_imag) - $signed(outputWires_2_real); // @[FixedPointTypeClass.scala 33:22]
  assign _GEN_2115 = {{1{outputWires_2_real[15]}},outputWires_2_real}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_396 = $signed(_GEN_2115) * $signed(_T_393); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2116 = {{1{twiddles_3_imag[15]}},twiddles_3_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_397 = $signed(_T_394) * $signed(_GEN_2116); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2117 = {{1{_GEN_135[15]}},_GEN_135}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_398 = $signed(_T_395) * $signed(_GEN_2117); // @[FixedPointTypeClass.scala 211:35]
  assign _T_399 = $signed(_T_396) - $signed(_T_397); // @[FixedPointTypeClass.scala 33:22]
  assign _T_400 = $signed(_T_396) + $signed(_T_398); // @[FixedPointTypeClass.scala 24:22]
  assign _T_406 = $signed(_T_399) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_407 = _T_406[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_410 = $signed(_T_400) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_411 = _T_410[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_418 = sdf_stages_4_io_cntr < 9'h10; // @[SDFChainRadix22.scala 328:32]
  assign _T_419 = sdf_stages_4_io_cntr < 9'h18; // @[SDFChainRadix22.scala 328:78]
  assign _T_420 = _T_419 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign _T_421 = _T_418 ? 1'h0 : _T_420; // @[SDFChainRadix22.scala 328:19]
  assign outputWires_3_real = sdf_stages_3_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _T_427 = 16'sh0 - $signed(outputWires_3_real); // @[FixedPointTypeClass.scala 39:43]
  assign outputWires_3_imag = sdf_stages_3_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _GEN_202 = 7'h21 == _T_201[6:0] ? 6'h2 : 6'h0; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_203 = 7'h22 == _T_201[6:0] ? 6'h4 : _GEN_202; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_204 = 7'h23 == _T_201[6:0] ? 6'h6 : _GEN_203; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_205 = 7'h24 == _T_201[6:0] ? 6'h8 : _GEN_204; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_206 = 7'h25 == _T_201[6:0] ? 6'ha : _GEN_205; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_207 = 7'h26 == _T_201[6:0] ? 6'hc : _GEN_206; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_208 = 7'h27 == _T_201[6:0] ? 6'he : _GEN_207; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_209 = 7'h28 == _T_201[6:0] ? 6'h10 : _GEN_208; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_210 = 7'h29 == _T_201[6:0] ? 6'h12 : _GEN_209; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_211 = 7'h2a == _T_201[6:0] ? 6'h14 : _GEN_210; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_212 = 7'h2b == _T_201[6:0] ? 6'h16 : _GEN_211; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_213 = 7'h2c == _T_201[6:0] ? 6'h18 : _GEN_212; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_214 = 7'h2d == _T_201[6:0] ? 6'h1a : _GEN_213; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_215 = 7'h2e == _T_201[6:0] ? 6'h1c : _GEN_214; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_216 = 7'h2f == _T_201[6:0] ? 6'h1e : _GEN_215; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_217 = 7'h30 == _T_201[6:0] ? 6'h20 : _GEN_216; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_218 = 7'h31 == _T_201[6:0] ? 6'h22 : _GEN_217; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_219 = 7'h32 == _T_201[6:0] ? 6'h23 : _GEN_218; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_220 = 7'h33 == _T_201[6:0] ? 6'h24 : _GEN_219; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_221 = 7'h34 == _T_201[6:0] ? 6'h26 : _GEN_220; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_222 = 7'h35 == _T_201[6:0] ? 6'h27 : _GEN_221; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_223 = 7'h36 == _T_201[6:0] ? 6'h28 : _GEN_222; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_224 = 7'h37 == _T_201[6:0] ? 6'h2a : _GEN_223; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_225 = 7'h38 == _T_201[6:0] ? 6'h2b : _GEN_224; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_226 = 7'h39 == _T_201[6:0] ? 6'h2c : _GEN_225; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_227 = 7'h3a == _T_201[6:0] ? 6'h2e : _GEN_226; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_228 = 7'h3b == _T_201[6:0] ? 6'h2f : _GEN_227; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_229 = 7'h3c == _T_201[6:0] ? 6'h30 : _GEN_228; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_230 = 7'h3d == _T_201[6:0] ? 6'h32 : _GEN_229; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_231 = 7'h3e == _T_201[6:0] ? 6'h33 : _GEN_230; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_232 = 7'h3f == _T_201[6:0] ? 6'h34 : _GEN_231; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_233 = 7'h40 == _T_201[6:0] ? 6'h0 : _GEN_232; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_234 = 7'h41 == _T_201[6:0] ? 6'h1 : _GEN_233; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_235 = 7'h42 == _T_201[6:0] ? 6'h2 : _GEN_234; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_236 = 7'h43 == _T_201[6:0] ? 6'h3 : _GEN_235; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_237 = 7'h44 == _T_201[6:0] ? 6'h4 : _GEN_236; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_238 = 7'h45 == _T_201[6:0] ? 6'h5 : _GEN_237; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_239 = 7'h46 == _T_201[6:0] ? 6'h6 : _GEN_238; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_240 = 7'h47 == _T_201[6:0] ? 6'h7 : _GEN_239; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_241 = 7'h48 == _T_201[6:0] ? 6'h8 : _GEN_240; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_242 = 7'h49 == _T_201[6:0] ? 6'h9 : _GEN_241; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_243 = 7'h4a == _T_201[6:0] ? 6'ha : _GEN_242; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_244 = 7'h4b == _T_201[6:0] ? 6'hb : _GEN_243; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_245 = 7'h4c == _T_201[6:0] ? 6'hc : _GEN_244; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_246 = 7'h4d == _T_201[6:0] ? 6'hd : _GEN_245; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_247 = 7'h4e == _T_201[6:0] ? 6'he : _GEN_246; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_248 = 7'h4f == _T_201[6:0] ? 6'hf : _GEN_247; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_249 = 7'h50 == _T_201[6:0] ? 6'h10 : _GEN_248; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_250 = 7'h51 == _T_201[6:0] ? 6'h11 : _GEN_249; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_251 = 7'h52 == _T_201[6:0] ? 6'h12 : _GEN_250; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_252 = 7'h53 == _T_201[6:0] ? 6'h13 : _GEN_251; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_253 = 7'h54 == _T_201[6:0] ? 6'h14 : _GEN_252; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_254 = 7'h55 == _T_201[6:0] ? 6'h15 : _GEN_253; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_255 = 7'h56 == _T_201[6:0] ? 6'h16 : _GEN_254; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_256 = 7'h57 == _T_201[6:0] ? 6'h17 : _GEN_255; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_257 = 7'h58 == _T_201[6:0] ? 6'h18 : _GEN_256; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_258 = 7'h59 == _T_201[6:0] ? 6'h19 : _GEN_257; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_259 = 7'h5a == _T_201[6:0] ? 6'h1a : _GEN_258; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_260 = 7'h5b == _T_201[6:0] ? 6'h1b : _GEN_259; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_261 = 7'h5c == _T_201[6:0] ? 6'h1c : _GEN_260; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_262 = 7'h5d == _T_201[6:0] ? 6'h1d : _GEN_261; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_263 = 7'h5e == _T_201[6:0] ? 6'h1e : _GEN_262; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_264 = 7'h5f == _T_201[6:0] ? 6'h1f : _GEN_263; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_265 = 7'h60 == _T_201[6:0] ? 6'h0 : _GEN_264; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_266 = 7'h61 == _T_201[6:0] ? 6'h3 : _GEN_265; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_267 = 7'h62 == _T_201[6:0] ? 6'h6 : _GEN_266; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_268 = 7'h63 == _T_201[6:0] ? 6'h9 : _GEN_267; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_269 = 7'h64 == _T_201[6:0] ? 6'hc : _GEN_268; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_270 = 7'h65 == _T_201[6:0] ? 6'hf : _GEN_269; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_271 = 7'h66 == _T_201[6:0] ? 6'h12 : _GEN_270; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_272 = 7'h67 == _T_201[6:0] ? 6'h15 : _GEN_271; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_273 = 7'h68 == _T_201[6:0] ? 6'h18 : _GEN_272; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_274 = 7'h69 == _T_201[6:0] ? 6'h1b : _GEN_273; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_275 = 7'h6a == _T_201[6:0] ? 6'h1e : _GEN_274; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_276 = 7'h6b == _T_201[6:0] ? 6'h21 : _GEN_275; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_277 = 7'h6c == _T_201[6:0] ? 6'h23 : _GEN_276; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_278 = 7'h6d == _T_201[6:0] ? 6'h25 : _GEN_277; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_279 = 7'h6e == _T_201[6:0] ? 6'h27 : _GEN_278; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_280 = 7'h6f == _T_201[6:0] ? 6'h29 : _GEN_279; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_281 = 7'h70 == _T_201[6:0] ? 6'h2b : _GEN_280; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_282 = 7'h71 == _T_201[6:0] ? 6'h2d : _GEN_281; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_283 = 7'h72 == _T_201[6:0] ? 6'h2f : _GEN_282; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_284 = 7'h73 == _T_201[6:0] ? 6'h31 : _GEN_283; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_285 = 7'h74 == _T_201[6:0] ? 6'h33 : _GEN_284; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_286 = 7'h75 == _T_201[6:0] ? 6'h35 : _GEN_285; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_287 = 7'h76 == _T_201[6:0] ? 6'h36 : _GEN_286; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_288 = 7'h77 == _T_201[6:0] ? 6'h37 : _GEN_287; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_289 = 7'h78 == _T_201[6:0] ? 6'h38 : _GEN_288; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_290 = 7'h79 == _T_201[6:0] ? 6'h39 : _GEN_289; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_291 = 7'h7a == _T_201[6:0] ? 6'h3a : _GEN_290; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_292 = 7'h7b == _T_201[6:0] ? 6'h3b : _GEN_291; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_293 = 7'h7c == _T_201[6:0] ? 6'h3c : _GEN_292; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_294 = 7'h7d == _T_201[6:0] ? 6'h3d : _GEN_293; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_295 = 7'h7e == _T_201[6:0] ? 6'h3e : _GEN_294; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_296 = 7'h7f == _T_201[6:0] ? 6'h3f : _GEN_295; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_299 = 6'h1 == _GEN_296 ? $signed(16'sh3fec) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_300 = 6'h1 == _GEN_296 ? $signed(-16'sh324) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_301 = 6'h2 == _GEN_296 ? $signed(16'sh3fb1) : $signed(_GEN_299); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_302 = 6'h2 == _GEN_296 ? $signed(-16'sh646) : $signed(_GEN_300); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_303 = 6'h3 == _GEN_296 ? $signed(16'sh3f4f) : $signed(_GEN_301); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_304 = 6'h3 == _GEN_296 ? $signed(-16'sh964) : $signed(_GEN_302); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_305 = 6'h4 == _GEN_296 ? $signed(16'sh3ec5) : $signed(_GEN_303); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_306 = 6'h4 == _GEN_296 ? $signed(-16'shc7c) : $signed(_GEN_304); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_307 = 6'h5 == _GEN_296 ? $signed(16'sh3e15) : $signed(_GEN_305); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_308 = 6'h5 == _GEN_296 ? $signed(-16'shf8d) : $signed(_GEN_306); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_309 = 6'h6 == _GEN_296 ? $signed(16'sh3d3f) : $signed(_GEN_307); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_310 = 6'h6 == _GEN_296 ? $signed(-16'sh1294) : $signed(_GEN_308); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_311 = 6'h7 == _GEN_296 ? $signed(16'sh3c42) : $signed(_GEN_309); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_312 = 6'h7 == _GEN_296 ? $signed(-16'sh1590) : $signed(_GEN_310); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_313 = 6'h8 == _GEN_296 ? $signed(16'sh3b21) : $signed(_GEN_311); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_314 = 6'h8 == _GEN_296 ? $signed(-16'sh187e) : $signed(_GEN_312); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_315 = 6'h9 == _GEN_296 ? $signed(16'sh39db) : $signed(_GEN_313); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_316 = 6'h9 == _GEN_296 ? $signed(-16'sh1b5d) : $signed(_GEN_314); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_317 = 6'ha == _GEN_296 ? $signed(16'sh3871) : $signed(_GEN_315); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_318 = 6'ha == _GEN_296 ? $signed(-16'sh1e2b) : $signed(_GEN_316); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_319 = 6'hb == _GEN_296 ? $signed(16'sh36e5) : $signed(_GEN_317); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_320 = 6'hb == _GEN_296 ? $signed(-16'sh20e7) : $signed(_GEN_318); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_321 = 6'hc == _GEN_296 ? $signed(16'sh3537) : $signed(_GEN_319); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_322 = 6'hc == _GEN_296 ? $signed(-16'sh238e) : $signed(_GEN_320); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_323 = 6'hd == _GEN_296 ? $signed(16'sh3368) : $signed(_GEN_321); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_324 = 6'hd == _GEN_296 ? $signed(-16'sh2620) : $signed(_GEN_322); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_325 = 6'he == _GEN_296 ? $signed(16'sh3179) : $signed(_GEN_323); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_326 = 6'he == _GEN_296 ? $signed(-16'sh289a) : $signed(_GEN_324); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_327 = 6'hf == _GEN_296 ? $signed(16'sh2f6c) : $signed(_GEN_325); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_328 = 6'hf == _GEN_296 ? $signed(-16'sh2afb) : $signed(_GEN_326); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_329 = 6'h10 == _GEN_296 ? $signed(16'sh2d41) : $signed(_GEN_327); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_330 = 6'h10 == _GEN_296 ? $signed(-16'sh2d41) : $signed(_GEN_328); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_331 = 6'h11 == _GEN_296 ? $signed(16'sh2afb) : $signed(_GEN_329); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_332 = 6'h11 == _GEN_296 ? $signed(-16'sh2f6c) : $signed(_GEN_330); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_333 = 6'h12 == _GEN_296 ? $signed(16'sh289a) : $signed(_GEN_331); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_334 = 6'h12 == _GEN_296 ? $signed(-16'sh3179) : $signed(_GEN_332); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_335 = 6'h13 == _GEN_296 ? $signed(16'sh2620) : $signed(_GEN_333); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_336 = 6'h13 == _GEN_296 ? $signed(-16'sh3368) : $signed(_GEN_334); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_337 = 6'h14 == _GEN_296 ? $signed(16'sh238e) : $signed(_GEN_335); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_338 = 6'h14 == _GEN_296 ? $signed(-16'sh3537) : $signed(_GEN_336); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_339 = 6'h15 == _GEN_296 ? $signed(16'sh20e7) : $signed(_GEN_337); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_340 = 6'h15 == _GEN_296 ? $signed(-16'sh36e5) : $signed(_GEN_338); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_341 = 6'h16 == _GEN_296 ? $signed(16'sh1e2b) : $signed(_GEN_339); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_342 = 6'h16 == _GEN_296 ? $signed(-16'sh3871) : $signed(_GEN_340); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_343 = 6'h17 == _GEN_296 ? $signed(16'sh1b5d) : $signed(_GEN_341); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_344 = 6'h17 == _GEN_296 ? $signed(-16'sh39db) : $signed(_GEN_342); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_345 = 6'h18 == _GEN_296 ? $signed(16'sh187e) : $signed(_GEN_343); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_346 = 6'h18 == _GEN_296 ? $signed(-16'sh3b21) : $signed(_GEN_344); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_347 = 6'h19 == _GEN_296 ? $signed(16'sh1590) : $signed(_GEN_345); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_348 = 6'h19 == _GEN_296 ? $signed(-16'sh3c42) : $signed(_GEN_346); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_349 = 6'h1a == _GEN_296 ? $signed(16'sh1294) : $signed(_GEN_347); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_350 = 6'h1a == _GEN_296 ? $signed(-16'sh3d3f) : $signed(_GEN_348); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_351 = 6'h1b == _GEN_296 ? $signed(16'shf8d) : $signed(_GEN_349); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_352 = 6'h1b == _GEN_296 ? $signed(-16'sh3e15) : $signed(_GEN_350); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_353 = 6'h1c == _GEN_296 ? $signed(16'shc7c) : $signed(_GEN_351); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_354 = 6'h1c == _GEN_296 ? $signed(-16'sh3ec5) : $signed(_GEN_352); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_355 = 6'h1d == _GEN_296 ? $signed(16'sh964) : $signed(_GEN_353); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_356 = 6'h1d == _GEN_296 ? $signed(-16'sh3f4f) : $signed(_GEN_354); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_357 = 6'h1e == _GEN_296 ? $signed(16'sh646) : $signed(_GEN_355); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_358 = 6'h1e == _GEN_296 ? $signed(-16'sh3fb1) : $signed(_GEN_356); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_359 = 6'h1f == _GEN_296 ? $signed(16'sh324) : $signed(_GEN_357); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_360 = 6'h1f == _GEN_296 ? $signed(-16'sh3fec) : $signed(_GEN_358); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_361 = 6'h20 == _GEN_296 ? $signed(16'sh0) : $signed(_GEN_359); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_362 = 6'h20 == _GEN_296 ? $signed(-16'sh4000) : $signed(_GEN_360); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_363 = 6'h21 == _GEN_296 ? $signed(-16'sh324) : $signed(_GEN_361); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_364 = 6'h21 == _GEN_296 ? $signed(-16'sh3fec) : $signed(_GEN_362); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_365 = 6'h22 == _GEN_296 ? $signed(-16'sh646) : $signed(_GEN_363); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_366 = 6'h22 == _GEN_296 ? $signed(-16'sh3fb1) : $signed(_GEN_364); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_367 = 6'h23 == _GEN_296 ? $signed(-16'shc7c) : $signed(_GEN_365); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_368 = 6'h23 == _GEN_296 ? $signed(-16'sh3ec5) : $signed(_GEN_366); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_369 = 6'h24 == _GEN_296 ? $signed(-16'sh1294) : $signed(_GEN_367); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_370 = 6'h24 == _GEN_296 ? $signed(-16'sh3d3f) : $signed(_GEN_368); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_371 = 6'h25 == _GEN_296 ? $signed(-16'sh1590) : $signed(_GEN_369); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_372 = 6'h25 == _GEN_296 ? $signed(-16'sh3c42) : $signed(_GEN_370); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_373 = 6'h26 == _GEN_296 ? $signed(-16'sh187e) : $signed(_GEN_371); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_374 = 6'h26 == _GEN_296 ? $signed(-16'sh3b21) : $signed(_GEN_372); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_375 = 6'h27 == _GEN_296 ? $signed(-16'sh1e2b) : $signed(_GEN_373); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_376 = 6'h27 == _GEN_296 ? $signed(-16'sh3871) : $signed(_GEN_374); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_377 = 6'h28 == _GEN_296 ? $signed(-16'sh238e) : $signed(_GEN_375); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_378 = 6'h28 == _GEN_296 ? $signed(-16'sh3537) : $signed(_GEN_376); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_379 = 6'h29 == _GEN_296 ? $signed(-16'sh2620) : $signed(_GEN_377); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_380 = 6'h29 == _GEN_296 ? $signed(-16'sh3368) : $signed(_GEN_378); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_381 = 6'h2a == _GEN_296 ? $signed(-16'sh289a) : $signed(_GEN_379); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_382 = 6'h2a == _GEN_296 ? $signed(-16'sh3179) : $signed(_GEN_380); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_383 = 6'h2b == _GEN_296 ? $signed(-16'sh2d41) : $signed(_GEN_381); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_384 = 6'h2b == _GEN_296 ? $signed(-16'sh2d41) : $signed(_GEN_382); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_385 = 6'h2c == _GEN_296 ? $signed(-16'sh3179) : $signed(_GEN_383); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_386 = 6'h2c == _GEN_296 ? $signed(-16'sh289a) : $signed(_GEN_384); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_387 = 6'h2d == _GEN_296 ? $signed(-16'sh3368) : $signed(_GEN_385); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_388 = 6'h2d == _GEN_296 ? $signed(-16'sh2620) : $signed(_GEN_386); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_389 = 6'h2e == _GEN_296 ? $signed(-16'sh3537) : $signed(_GEN_387); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_390 = 6'h2e == _GEN_296 ? $signed(-16'sh238e) : $signed(_GEN_388); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_391 = 6'h2f == _GEN_296 ? $signed(-16'sh3871) : $signed(_GEN_389); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_392 = 6'h2f == _GEN_296 ? $signed(-16'sh1e2b) : $signed(_GEN_390); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_393 = 6'h30 == _GEN_296 ? $signed(-16'sh3b21) : $signed(_GEN_391); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_394 = 6'h30 == _GEN_296 ? $signed(-16'sh187e) : $signed(_GEN_392); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_395 = 6'h31 == _GEN_296 ? $signed(-16'sh3c42) : $signed(_GEN_393); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_396 = 6'h31 == _GEN_296 ? $signed(-16'sh1590) : $signed(_GEN_394); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_397 = 6'h32 == _GEN_296 ? $signed(-16'sh3d3f) : $signed(_GEN_395); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_398 = 6'h32 == _GEN_296 ? $signed(-16'sh1294) : $signed(_GEN_396); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_399 = 6'h33 == _GEN_296 ? $signed(-16'sh3ec5) : $signed(_GEN_397); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_400 = 6'h33 == _GEN_296 ? $signed(-16'shc7c) : $signed(_GEN_398); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_401 = 6'h34 == _GEN_296 ? $signed(-16'sh3fb1) : $signed(_GEN_399); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_402 = 6'h34 == _GEN_296 ? $signed(-16'sh646) : $signed(_GEN_400); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_403 = 6'h35 == _GEN_296 ? $signed(-16'sh3fec) : $signed(_GEN_401); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_404 = 6'h35 == _GEN_296 ? $signed(-16'sh324) : $signed(_GEN_402); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_405 = 6'h36 == _GEN_296 ? $signed(-16'sh3fb1) : $signed(_GEN_403); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_406 = 6'h36 == _GEN_296 ? $signed(16'sh646) : $signed(_GEN_404); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_407 = 6'h37 == _GEN_296 ? $signed(-16'sh3e15) : $signed(_GEN_405); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_408 = 6'h37 == _GEN_296 ? $signed(16'shf8d) : $signed(_GEN_406); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_409 = 6'h38 == _GEN_296 ? $signed(-16'sh3b21) : $signed(_GEN_407); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_410 = 6'h38 == _GEN_296 ? $signed(16'sh187e) : $signed(_GEN_408); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_411 = 6'h39 == _GEN_296 ? $signed(-16'sh36e5) : $signed(_GEN_409); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_412 = 6'h39 == _GEN_296 ? $signed(16'sh20e7) : $signed(_GEN_410); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_413 = 6'h3a == _GEN_296 ? $signed(-16'sh3179) : $signed(_GEN_411); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_414 = 6'h3a == _GEN_296 ? $signed(16'sh289a) : $signed(_GEN_412); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_415 = 6'h3b == _GEN_296 ? $signed(-16'sh2afb) : $signed(_GEN_413); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_416 = 6'h3b == _GEN_296 ? $signed(16'sh2f6c) : $signed(_GEN_414); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_417 = 6'h3c == _GEN_296 ? $signed(-16'sh238e) : $signed(_GEN_415); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_418 = 6'h3c == _GEN_296 ? $signed(16'sh3537) : $signed(_GEN_416); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_419 = 6'h3d == _GEN_296 ? $signed(-16'sh1b5d) : $signed(_GEN_417); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_420 = 6'h3d == _GEN_296 ? $signed(16'sh39db) : $signed(_GEN_418); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_421 = 6'h3e == _GEN_296 ? $signed(-16'sh1294) : $signed(_GEN_419); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_422 = 6'h3e == _GEN_296 ? $signed(16'sh3d3f) : $signed(_GEN_420); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_423 = 6'h3f == _GEN_296 ? $signed(-16'sh964) : $signed(_GEN_421); // @[SDFChainRadix22.scala 291:27]
  assign twiddles_5_imag = 6'h3f == _GEN_296 ? $signed(16'sh3f4f) : $signed(_GEN_422); // @[SDFChainRadix22.scala 291:27]
  assign _T_765 = $signed(_GEN_423) + $signed(twiddles_5_imag); // @[FixedPointTypeClass.scala 24:22]
  assign outputWires_4_real = sdf_stages_4_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign outputWires_4_imag = sdf_stages_4_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign _T_766 = $signed(outputWires_4_real) + $signed(outputWires_4_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_767 = $signed(outputWires_4_imag) - $signed(outputWires_4_real); // @[FixedPointTypeClass.scala 33:22]
  assign _GEN_2118 = {{1{outputWires_4_real[15]}},outputWires_4_real}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_768 = $signed(_GEN_2118) * $signed(_T_765); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2119 = {{1{twiddles_5_imag[15]}},twiddles_5_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_769 = $signed(_T_766) * $signed(_GEN_2119); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2120 = {{1{_GEN_423[15]}},_GEN_423}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_770 = $signed(_T_767) * $signed(_GEN_2120); // @[FixedPointTypeClass.scala 211:35]
  assign _T_771 = $signed(_T_768) - $signed(_T_769); // @[FixedPointTypeClass.scala 33:22]
  assign _T_772 = $signed(_T_768) + $signed(_T_770); // @[FixedPointTypeClass.scala 24:22]
  assign _T_778 = $signed(_T_771) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_779 = _T_778[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_782 = $signed(_T_772) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_783 = _T_782[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_790 = sdf_stages_6_io_cntr < 9'h40; // @[SDFChainRadix22.scala 328:32]
  assign _T_791 = sdf_stages_6_io_cntr < 9'h60; // @[SDFChainRadix22.scala 328:78]
  assign _T_792 = _T_791 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign _T_793 = _T_790 ? 1'h0 : _T_792; // @[SDFChainRadix22.scala 328:19]
  assign outputWires_5_real = sdf_stages_5_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _T_799 = 16'sh0 - $signed(outputWires_5_real); // @[FixedPointTypeClass.scala 39:43]
  assign outputWires_5_imag = sdf_stages_5_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _GEN_682 = 9'h81 == _T_215 ? 8'h2 : 8'h0; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_683 = 9'h82 == _T_215 ? 8'h4 : _GEN_682; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_684 = 9'h83 == _T_215 ? 8'h6 : _GEN_683; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_685 = 9'h84 == _T_215 ? 8'h8 : _GEN_684; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_686 = 9'h85 == _T_215 ? 8'ha : _GEN_685; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_687 = 9'h86 == _T_215 ? 8'hc : _GEN_686; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_688 = 9'h87 == _T_215 ? 8'he : _GEN_687; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_689 = 9'h88 == _T_215 ? 8'h10 : _GEN_688; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_690 = 9'h89 == _T_215 ? 8'h12 : _GEN_689; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_691 = 9'h8a == _T_215 ? 8'h14 : _GEN_690; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_692 = 9'h8b == _T_215 ? 8'h16 : _GEN_691; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_693 = 9'h8c == _T_215 ? 8'h18 : _GEN_692; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_694 = 9'h8d == _T_215 ? 8'h1a : _GEN_693; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_695 = 9'h8e == _T_215 ? 8'h1c : _GEN_694; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_696 = 9'h8f == _T_215 ? 8'h1e : _GEN_695; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_697 = 9'h90 == _T_215 ? 8'h20 : _GEN_696; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_698 = 9'h91 == _T_215 ? 8'h22 : _GEN_697; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_699 = 9'h92 == _T_215 ? 8'h24 : _GEN_698; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_700 = 9'h93 == _T_215 ? 8'h26 : _GEN_699; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_701 = 9'h94 == _T_215 ? 8'h28 : _GEN_700; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_702 = 9'h95 == _T_215 ? 8'h2a : _GEN_701; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_703 = 9'h96 == _T_215 ? 8'h2c : _GEN_702; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_704 = 9'h97 == _T_215 ? 8'h2e : _GEN_703; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_705 = 9'h98 == _T_215 ? 8'h30 : _GEN_704; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_706 = 9'h99 == _T_215 ? 8'h32 : _GEN_705; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_707 = 9'h9a == _T_215 ? 8'h34 : _GEN_706; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_708 = 9'h9b == _T_215 ? 8'h36 : _GEN_707; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_709 = 9'h9c == _T_215 ? 8'h38 : _GEN_708; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_710 = 9'h9d == _T_215 ? 8'h3a : _GEN_709; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_711 = 9'h9e == _T_215 ? 8'h3c : _GEN_710; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_712 = 9'h9f == _T_215 ? 8'h3e : _GEN_711; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_713 = 9'ha0 == _T_215 ? 8'h40 : _GEN_712; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_714 = 9'ha1 == _T_215 ? 8'h42 : _GEN_713; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_715 = 9'ha2 == _T_215 ? 8'h44 : _GEN_714; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_716 = 9'ha3 == _T_215 ? 8'h46 : _GEN_715; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_717 = 9'ha4 == _T_215 ? 8'h48 : _GEN_716; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_718 = 9'ha5 == _T_215 ? 8'h4a : _GEN_717; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_719 = 9'ha6 == _T_215 ? 8'h4c : _GEN_718; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_720 = 9'ha7 == _T_215 ? 8'h4e : _GEN_719; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_721 = 9'ha8 == _T_215 ? 8'h50 : _GEN_720; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_722 = 9'ha9 == _T_215 ? 8'h52 : _GEN_721; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_723 = 9'haa == _T_215 ? 8'h54 : _GEN_722; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_724 = 9'hab == _T_215 ? 8'h56 : _GEN_723; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_725 = 9'hac == _T_215 ? 8'h58 : _GEN_724; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_726 = 9'had == _T_215 ? 8'h5a : _GEN_725; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_727 = 9'hae == _T_215 ? 8'h5c : _GEN_726; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_728 = 9'haf == _T_215 ? 8'h5e : _GEN_727; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_729 = 9'hb0 == _T_215 ? 8'h60 : _GEN_728; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_730 = 9'hb1 == _T_215 ? 8'h62 : _GEN_729; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_731 = 9'hb2 == _T_215 ? 8'h64 : _GEN_730; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_732 = 9'hb3 == _T_215 ? 8'h66 : _GEN_731; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_733 = 9'hb4 == _T_215 ? 8'h68 : _GEN_732; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_734 = 9'hb5 == _T_215 ? 8'h6a : _GEN_733; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_735 = 9'hb6 == _T_215 ? 8'h6c : _GEN_734; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_736 = 9'hb7 == _T_215 ? 8'h6e : _GEN_735; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_737 = 9'hb8 == _T_215 ? 8'h70 : _GEN_736; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_738 = 9'hb9 == _T_215 ? 8'h72 : _GEN_737; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_739 = 9'hba == _T_215 ? 8'h74 : _GEN_738; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_740 = 9'hbb == _T_215 ? 8'h76 : _GEN_739; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_741 = 9'hbc == _T_215 ? 8'h78 : _GEN_740; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_742 = 9'hbd == _T_215 ? 8'h7a : _GEN_741; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_743 = 9'hbe == _T_215 ? 8'h7c : _GEN_742; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_744 = 9'hbf == _T_215 ? 8'h7e : _GEN_743; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_745 = 9'hc0 == _T_215 ? 8'h80 : _GEN_744; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_746 = 9'hc1 == _T_215 ? 8'h82 : _GEN_745; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_747 = 9'hc2 == _T_215 ? 8'h83 : _GEN_746; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_748 = 9'hc3 == _T_215 ? 8'h84 : _GEN_747; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_749 = 9'hc4 == _T_215 ? 8'h86 : _GEN_748; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_750 = 9'hc5 == _T_215 ? 8'h87 : _GEN_749; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_751 = 9'hc6 == _T_215 ? 8'h88 : _GEN_750; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_752 = 9'hc7 == _T_215 ? 8'h8a : _GEN_751; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_753 = 9'hc8 == _T_215 ? 8'h8b : _GEN_752; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_754 = 9'hc9 == _T_215 ? 8'h8c : _GEN_753; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_755 = 9'hca == _T_215 ? 8'h8e : _GEN_754; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_756 = 9'hcb == _T_215 ? 8'h8f : _GEN_755; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_757 = 9'hcc == _T_215 ? 8'h90 : _GEN_756; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_758 = 9'hcd == _T_215 ? 8'h92 : _GEN_757; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_759 = 9'hce == _T_215 ? 8'h93 : _GEN_758; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_760 = 9'hcf == _T_215 ? 8'h94 : _GEN_759; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_761 = 9'hd0 == _T_215 ? 8'h96 : _GEN_760; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_762 = 9'hd1 == _T_215 ? 8'h97 : _GEN_761; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_763 = 9'hd2 == _T_215 ? 8'h98 : _GEN_762; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_764 = 9'hd3 == _T_215 ? 8'h9a : _GEN_763; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_765 = 9'hd4 == _T_215 ? 8'h9b : _GEN_764; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_766 = 9'hd5 == _T_215 ? 8'h9c : _GEN_765; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_767 = 9'hd6 == _T_215 ? 8'h9e : _GEN_766; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_768 = 9'hd7 == _T_215 ? 8'h9f : _GEN_767; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_769 = 9'hd8 == _T_215 ? 8'ha0 : _GEN_768; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_770 = 9'hd9 == _T_215 ? 8'ha2 : _GEN_769; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_771 = 9'hda == _T_215 ? 8'ha3 : _GEN_770; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_772 = 9'hdb == _T_215 ? 8'ha4 : _GEN_771; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_773 = 9'hdc == _T_215 ? 8'ha6 : _GEN_772; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_774 = 9'hdd == _T_215 ? 8'ha7 : _GEN_773; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_775 = 9'hde == _T_215 ? 8'ha8 : _GEN_774; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_776 = 9'hdf == _T_215 ? 8'haa : _GEN_775; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_777 = 9'he0 == _T_215 ? 8'hab : _GEN_776; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_778 = 9'he1 == _T_215 ? 8'hac : _GEN_777; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_779 = 9'he2 == _T_215 ? 8'hae : _GEN_778; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_780 = 9'he3 == _T_215 ? 8'haf : _GEN_779; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_781 = 9'he4 == _T_215 ? 8'hb0 : _GEN_780; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_782 = 9'he5 == _T_215 ? 8'hb2 : _GEN_781; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_783 = 9'he6 == _T_215 ? 8'hb3 : _GEN_782; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_784 = 9'he7 == _T_215 ? 8'hb4 : _GEN_783; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_785 = 9'he8 == _T_215 ? 8'hb6 : _GEN_784; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_786 = 9'he9 == _T_215 ? 8'hb7 : _GEN_785; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_787 = 9'hea == _T_215 ? 8'hb8 : _GEN_786; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_788 = 9'heb == _T_215 ? 8'hba : _GEN_787; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_789 = 9'hec == _T_215 ? 8'hbb : _GEN_788; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_790 = 9'hed == _T_215 ? 8'hbc : _GEN_789; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_791 = 9'hee == _T_215 ? 8'hbe : _GEN_790; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_792 = 9'hef == _T_215 ? 8'hbf : _GEN_791; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_793 = 9'hf0 == _T_215 ? 8'hc0 : _GEN_792; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_794 = 9'hf1 == _T_215 ? 8'hc2 : _GEN_793; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_795 = 9'hf2 == _T_215 ? 8'hc3 : _GEN_794; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_796 = 9'hf3 == _T_215 ? 8'hc4 : _GEN_795; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_797 = 9'hf4 == _T_215 ? 8'hc6 : _GEN_796; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_798 = 9'hf5 == _T_215 ? 8'hc7 : _GEN_797; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_799 = 9'hf6 == _T_215 ? 8'hc8 : _GEN_798; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_800 = 9'hf7 == _T_215 ? 8'hca : _GEN_799; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_801 = 9'hf8 == _T_215 ? 8'hcb : _GEN_800; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_802 = 9'hf9 == _T_215 ? 8'hcc : _GEN_801; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_803 = 9'hfa == _T_215 ? 8'hce : _GEN_802; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_804 = 9'hfb == _T_215 ? 8'hcf : _GEN_803; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_805 = 9'hfc == _T_215 ? 8'hd0 : _GEN_804; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_806 = 9'hfd == _T_215 ? 8'hd2 : _GEN_805; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_807 = 9'hfe == _T_215 ? 8'hd3 : _GEN_806; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_808 = 9'hff == _T_215 ? 8'hd4 : _GEN_807; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_809 = 9'h100 == _T_215 ? 8'h0 : _GEN_808; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_810 = 9'h101 == _T_215 ? 8'h1 : _GEN_809; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_811 = 9'h102 == _T_215 ? 8'h2 : _GEN_810; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_812 = 9'h103 == _T_215 ? 8'h3 : _GEN_811; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_813 = 9'h104 == _T_215 ? 8'h4 : _GEN_812; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_814 = 9'h105 == _T_215 ? 8'h5 : _GEN_813; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_815 = 9'h106 == _T_215 ? 8'h6 : _GEN_814; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_816 = 9'h107 == _T_215 ? 8'h7 : _GEN_815; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_817 = 9'h108 == _T_215 ? 8'h8 : _GEN_816; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_818 = 9'h109 == _T_215 ? 8'h9 : _GEN_817; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_819 = 9'h10a == _T_215 ? 8'ha : _GEN_818; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_820 = 9'h10b == _T_215 ? 8'hb : _GEN_819; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_821 = 9'h10c == _T_215 ? 8'hc : _GEN_820; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_822 = 9'h10d == _T_215 ? 8'hd : _GEN_821; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_823 = 9'h10e == _T_215 ? 8'he : _GEN_822; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_824 = 9'h10f == _T_215 ? 8'hf : _GEN_823; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_825 = 9'h110 == _T_215 ? 8'h10 : _GEN_824; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_826 = 9'h111 == _T_215 ? 8'h11 : _GEN_825; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_827 = 9'h112 == _T_215 ? 8'h12 : _GEN_826; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_828 = 9'h113 == _T_215 ? 8'h13 : _GEN_827; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_829 = 9'h114 == _T_215 ? 8'h14 : _GEN_828; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_830 = 9'h115 == _T_215 ? 8'h15 : _GEN_829; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_831 = 9'h116 == _T_215 ? 8'h16 : _GEN_830; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_832 = 9'h117 == _T_215 ? 8'h17 : _GEN_831; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_833 = 9'h118 == _T_215 ? 8'h18 : _GEN_832; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_834 = 9'h119 == _T_215 ? 8'h19 : _GEN_833; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_835 = 9'h11a == _T_215 ? 8'h1a : _GEN_834; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_836 = 9'h11b == _T_215 ? 8'h1b : _GEN_835; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_837 = 9'h11c == _T_215 ? 8'h1c : _GEN_836; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_838 = 9'h11d == _T_215 ? 8'h1d : _GEN_837; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_839 = 9'h11e == _T_215 ? 8'h1e : _GEN_838; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_840 = 9'h11f == _T_215 ? 8'h1f : _GEN_839; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_841 = 9'h120 == _T_215 ? 8'h20 : _GEN_840; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_842 = 9'h121 == _T_215 ? 8'h21 : _GEN_841; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_843 = 9'h122 == _T_215 ? 8'h22 : _GEN_842; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_844 = 9'h123 == _T_215 ? 8'h23 : _GEN_843; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_845 = 9'h124 == _T_215 ? 8'h24 : _GEN_844; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_846 = 9'h125 == _T_215 ? 8'h25 : _GEN_845; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_847 = 9'h126 == _T_215 ? 8'h26 : _GEN_846; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_848 = 9'h127 == _T_215 ? 8'h27 : _GEN_847; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_849 = 9'h128 == _T_215 ? 8'h28 : _GEN_848; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_850 = 9'h129 == _T_215 ? 8'h29 : _GEN_849; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_851 = 9'h12a == _T_215 ? 8'h2a : _GEN_850; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_852 = 9'h12b == _T_215 ? 8'h2b : _GEN_851; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_853 = 9'h12c == _T_215 ? 8'h2c : _GEN_852; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_854 = 9'h12d == _T_215 ? 8'h2d : _GEN_853; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_855 = 9'h12e == _T_215 ? 8'h2e : _GEN_854; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_856 = 9'h12f == _T_215 ? 8'h2f : _GEN_855; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_857 = 9'h130 == _T_215 ? 8'h30 : _GEN_856; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_858 = 9'h131 == _T_215 ? 8'h31 : _GEN_857; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_859 = 9'h132 == _T_215 ? 8'h32 : _GEN_858; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_860 = 9'h133 == _T_215 ? 8'h33 : _GEN_859; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_861 = 9'h134 == _T_215 ? 8'h34 : _GEN_860; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_862 = 9'h135 == _T_215 ? 8'h35 : _GEN_861; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_863 = 9'h136 == _T_215 ? 8'h36 : _GEN_862; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_864 = 9'h137 == _T_215 ? 8'h37 : _GEN_863; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_865 = 9'h138 == _T_215 ? 8'h38 : _GEN_864; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_866 = 9'h139 == _T_215 ? 8'h39 : _GEN_865; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_867 = 9'h13a == _T_215 ? 8'h3a : _GEN_866; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_868 = 9'h13b == _T_215 ? 8'h3b : _GEN_867; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_869 = 9'h13c == _T_215 ? 8'h3c : _GEN_868; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_870 = 9'h13d == _T_215 ? 8'h3d : _GEN_869; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_871 = 9'h13e == _T_215 ? 8'h3e : _GEN_870; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_872 = 9'h13f == _T_215 ? 8'h3f : _GEN_871; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_873 = 9'h140 == _T_215 ? 8'h40 : _GEN_872; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_874 = 9'h141 == _T_215 ? 8'h41 : _GEN_873; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_875 = 9'h142 == _T_215 ? 8'h42 : _GEN_874; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_876 = 9'h143 == _T_215 ? 8'h43 : _GEN_875; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_877 = 9'h144 == _T_215 ? 8'h44 : _GEN_876; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_878 = 9'h145 == _T_215 ? 8'h45 : _GEN_877; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_879 = 9'h146 == _T_215 ? 8'h46 : _GEN_878; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_880 = 9'h147 == _T_215 ? 8'h47 : _GEN_879; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_881 = 9'h148 == _T_215 ? 8'h48 : _GEN_880; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_882 = 9'h149 == _T_215 ? 8'h49 : _GEN_881; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_883 = 9'h14a == _T_215 ? 8'h4a : _GEN_882; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_884 = 9'h14b == _T_215 ? 8'h4b : _GEN_883; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_885 = 9'h14c == _T_215 ? 8'h4c : _GEN_884; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_886 = 9'h14d == _T_215 ? 8'h4d : _GEN_885; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_887 = 9'h14e == _T_215 ? 8'h4e : _GEN_886; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_888 = 9'h14f == _T_215 ? 8'h4f : _GEN_887; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_889 = 9'h150 == _T_215 ? 8'h50 : _GEN_888; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_890 = 9'h151 == _T_215 ? 8'h51 : _GEN_889; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_891 = 9'h152 == _T_215 ? 8'h52 : _GEN_890; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_892 = 9'h153 == _T_215 ? 8'h53 : _GEN_891; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_893 = 9'h154 == _T_215 ? 8'h54 : _GEN_892; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_894 = 9'h155 == _T_215 ? 8'h55 : _GEN_893; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_895 = 9'h156 == _T_215 ? 8'h56 : _GEN_894; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_896 = 9'h157 == _T_215 ? 8'h57 : _GEN_895; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_897 = 9'h158 == _T_215 ? 8'h58 : _GEN_896; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_898 = 9'h159 == _T_215 ? 8'h59 : _GEN_897; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_899 = 9'h15a == _T_215 ? 8'h5a : _GEN_898; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_900 = 9'h15b == _T_215 ? 8'h5b : _GEN_899; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_901 = 9'h15c == _T_215 ? 8'h5c : _GEN_900; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_902 = 9'h15d == _T_215 ? 8'h5d : _GEN_901; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_903 = 9'h15e == _T_215 ? 8'h5e : _GEN_902; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_904 = 9'h15f == _T_215 ? 8'h5f : _GEN_903; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_905 = 9'h160 == _T_215 ? 8'h60 : _GEN_904; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_906 = 9'h161 == _T_215 ? 8'h61 : _GEN_905; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_907 = 9'h162 == _T_215 ? 8'h62 : _GEN_906; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_908 = 9'h163 == _T_215 ? 8'h63 : _GEN_907; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_909 = 9'h164 == _T_215 ? 8'h64 : _GEN_908; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_910 = 9'h165 == _T_215 ? 8'h65 : _GEN_909; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_911 = 9'h166 == _T_215 ? 8'h66 : _GEN_910; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_912 = 9'h167 == _T_215 ? 8'h67 : _GEN_911; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_913 = 9'h168 == _T_215 ? 8'h68 : _GEN_912; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_914 = 9'h169 == _T_215 ? 8'h69 : _GEN_913; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_915 = 9'h16a == _T_215 ? 8'h6a : _GEN_914; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_916 = 9'h16b == _T_215 ? 8'h6b : _GEN_915; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_917 = 9'h16c == _T_215 ? 8'h6c : _GEN_916; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_918 = 9'h16d == _T_215 ? 8'h6d : _GEN_917; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_919 = 9'h16e == _T_215 ? 8'h6e : _GEN_918; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_920 = 9'h16f == _T_215 ? 8'h6f : _GEN_919; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_921 = 9'h170 == _T_215 ? 8'h70 : _GEN_920; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_922 = 9'h171 == _T_215 ? 8'h71 : _GEN_921; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_923 = 9'h172 == _T_215 ? 8'h72 : _GEN_922; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_924 = 9'h173 == _T_215 ? 8'h73 : _GEN_923; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_925 = 9'h174 == _T_215 ? 8'h74 : _GEN_924; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_926 = 9'h175 == _T_215 ? 8'h75 : _GEN_925; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_927 = 9'h176 == _T_215 ? 8'h76 : _GEN_926; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_928 = 9'h177 == _T_215 ? 8'h77 : _GEN_927; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_929 = 9'h178 == _T_215 ? 8'h78 : _GEN_928; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_930 = 9'h179 == _T_215 ? 8'h79 : _GEN_929; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_931 = 9'h17a == _T_215 ? 8'h7a : _GEN_930; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_932 = 9'h17b == _T_215 ? 8'h7b : _GEN_931; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_933 = 9'h17c == _T_215 ? 8'h7c : _GEN_932; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_934 = 9'h17d == _T_215 ? 8'h7d : _GEN_933; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_935 = 9'h17e == _T_215 ? 8'h7e : _GEN_934; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_936 = 9'h17f == _T_215 ? 8'h7f : _GEN_935; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_937 = 9'h180 == _T_215 ? 8'h0 : _GEN_936; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_938 = 9'h181 == _T_215 ? 8'h3 : _GEN_937; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_939 = 9'h182 == _T_215 ? 8'h6 : _GEN_938; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_940 = 9'h183 == _T_215 ? 8'h9 : _GEN_939; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_941 = 9'h184 == _T_215 ? 8'hc : _GEN_940; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_942 = 9'h185 == _T_215 ? 8'hf : _GEN_941; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_943 = 9'h186 == _T_215 ? 8'h12 : _GEN_942; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_944 = 9'h187 == _T_215 ? 8'h15 : _GEN_943; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_945 = 9'h188 == _T_215 ? 8'h18 : _GEN_944; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_946 = 9'h189 == _T_215 ? 8'h1b : _GEN_945; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_947 = 9'h18a == _T_215 ? 8'h1e : _GEN_946; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_948 = 9'h18b == _T_215 ? 8'h21 : _GEN_947; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_949 = 9'h18c == _T_215 ? 8'h24 : _GEN_948; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_950 = 9'h18d == _T_215 ? 8'h27 : _GEN_949; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_951 = 9'h18e == _T_215 ? 8'h2a : _GEN_950; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_952 = 9'h18f == _T_215 ? 8'h2d : _GEN_951; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_953 = 9'h190 == _T_215 ? 8'h30 : _GEN_952; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_954 = 9'h191 == _T_215 ? 8'h33 : _GEN_953; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_955 = 9'h192 == _T_215 ? 8'h36 : _GEN_954; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_956 = 9'h193 == _T_215 ? 8'h39 : _GEN_955; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_957 = 9'h194 == _T_215 ? 8'h3c : _GEN_956; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_958 = 9'h195 == _T_215 ? 8'h3f : _GEN_957; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_959 = 9'h196 == _T_215 ? 8'h42 : _GEN_958; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_960 = 9'h197 == _T_215 ? 8'h45 : _GEN_959; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_961 = 9'h198 == _T_215 ? 8'h48 : _GEN_960; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_962 = 9'h199 == _T_215 ? 8'h4b : _GEN_961; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_963 = 9'h19a == _T_215 ? 8'h4e : _GEN_962; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_964 = 9'h19b == _T_215 ? 8'h51 : _GEN_963; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_965 = 9'h19c == _T_215 ? 8'h54 : _GEN_964; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_966 = 9'h19d == _T_215 ? 8'h57 : _GEN_965; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_967 = 9'h19e == _T_215 ? 8'h5a : _GEN_966; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_968 = 9'h19f == _T_215 ? 8'h5d : _GEN_967; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_969 = 9'h1a0 == _T_215 ? 8'h60 : _GEN_968; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_970 = 9'h1a1 == _T_215 ? 8'h63 : _GEN_969; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_971 = 9'h1a2 == _T_215 ? 8'h66 : _GEN_970; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_972 = 9'h1a3 == _T_215 ? 8'h69 : _GEN_971; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_973 = 9'h1a4 == _T_215 ? 8'h6c : _GEN_972; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_974 = 9'h1a5 == _T_215 ? 8'h6f : _GEN_973; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_975 = 9'h1a6 == _T_215 ? 8'h72 : _GEN_974; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_976 = 9'h1a7 == _T_215 ? 8'h75 : _GEN_975; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_977 = 9'h1a8 == _T_215 ? 8'h78 : _GEN_976; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_978 = 9'h1a9 == _T_215 ? 8'h7b : _GEN_977; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_979 = 9'h1aa == _T_215 ? 8'h7e : _GEN_978; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_980 = 9'h1ab == _T_215 ? 8'h81 : _GEN_979; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_981 = 9'h1ac == _T_215 ? 8'h83 : _GEN_980; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_982 = 9'h1ad == _T_215 ? 8'h85 : _GEN_981; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_983 = 9'h1ae == _T_215 ? 8'h87 : _GEN_982; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_984 = 9'h1af == _T_215 ? 8'h89 : _GEN_983; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_985 = 9'h1b0 == _T_215 ? 8'h8b : _GEN_984; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_986 = 9'h1b1 == _T_215 ? 8'h8d : _GEN_985; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_987 = 9'h1b2 == _T_215 ? 8'h8f : _GEN_986; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_988 = 9'h1b3 == _T_215 ? 8'h91 : _GEN_987; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_989 = 9'h1b4 == _T_215 ? 8'h93 : _GEN_988; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_990 = 9'h1b5 == _T_215 ? 8'h95 : _GEN_989; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_991 = 9'h1b6 == _T_215 ? 8'h97 : _GEN_990; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_992 = 9'h1b7 == _T_215 ? 8'h99 : _GEN_991; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_993 = 9'h1b8 == _T_215 ? 8'h9b : _GEN_992; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_994 = 9'h1b9 == _T_215 ? 8'h9d : _GEN_993; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_995 = 9'h1ba == _T_215 ? 8'h9f : _GEN_994; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_996 = 9'h1bb == _T_215 ? 8'ha1 : _GEN_995; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_997 = 9'h1bc == _T_215 ? 8'ha3 : _GEN_996; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_998 = 9'h1bd == _T_215 ? 8'ha5 : _GEN_997; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_999 = 9'h1be == _T_215 ? 8'ha7 : _GEN_998; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1000 = 9'h1bf == _T_215 ? 8'ha9 : _GEN_999; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1001 = 9'h1c0 == _T_215 ? 8'hab : _GEN_1000; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1002 = 9'h1c1 == _T_215 ? 8'had : _GEN_1001; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1003 = 9'h1c2 == _T_215 ? 8'haf : _GEN_1002; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1004 = 9'h1c3 == _T_215 ? 8'hb1 : _GEN_1003; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1005 = 9'h1c4 == _T_215 ? 8'hb3 : _GEN_1004; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1006 = 9'h1c5 == _T_215 ? 8'hb5 : _GEN_1005; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1007 = 9'h1c6 == _T_215 ? 8'hb7 : _GEN_1006; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1008 = 9'h1c7 == _T_215 ? 8'hb9 : _GEN_1007; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1009 = 9'h1c8 == _T_215 ? 8'hbb : _GEN_1008; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1010 = 9'h1c9 == _T_215 ? 8'hbd : _GEN_1009; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1011 = 9'h1ca == _T_215 ? 8'hbf : _GEN_1010; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1012 = 9'h1cb == _T_215 ? 8'hc1 : _GEN_1011; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1013 = 9'h1cc == _T_215 ? 8'hc3 : _GEN_1012; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1014 = 9'h1cd == _T_215 ? 8'hc5 : _GEN_1013; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1015 = 9'h1ce == _T_215 ? 8'hc7 : _GEN_1014; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1016 = 9'h1cf == _T_215 ? 8'hc9 : _GEN_1015; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1017 = 9'h1d0 == _T_215 ? 8'hcb : _GEN_1016; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1018 = 9'h1d1 == _T_215 ? 8'hcd : _GEN_1017; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1019 = 9'h1d2 == _T_215 ? 8'hcf : _GEN_1018; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1020 = 9'h1d3 == _T_215 ? 8'hd1 : _GEN_1019; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1021 = 9'h1d4 == _T_215 ? 8'hd3 : _GEN_1020; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1022 = 9'h1d5 == _T_215 ? 8'hd5 : _GEN_1021; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1023 = 9'h1d6 == _T_215 ? 8'hd6 : _GEN_1022; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1024 = 9'h1d7 == _T_215 ? 8'hd7 : _GEN_1023; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1025 = 9'h1d8 == _T_215 ? 8'hd8 : _GEN_1024; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1026 = 9'h1d9 == _T_215 ? 8'hd9 : _GEN_1025; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1027 = 9'h1da == _T_215 ? 8'hda : _GEN_1026; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1028 = 9'h1db == _T_215 ? 8'hdb : _GEN_1027; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1029 = 9'h1dc == _T_215 ? 8'hdc : _GEN_1028; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1030 = 9'h1dd == _T_215 ? 8'hdd : _GEN_1029; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1031 = 9'h1de == _T_215 ? 8'hde : _GEN_1030; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1032 = 9'h1df == _T_215 ? 8'hdf : _GEN_1031; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1033 = 9'h1e0 == _T_215 ? 8'he0 : _GEN_1032; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1034 = 9'h1e1 == _T_215 ? 8'he1 : _GEN_1033; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1035 = 9'h1e2 == _T_215 ? 8'he2 : _GEN_1034; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1036 = 9'h1e3 == _T_215 ? 8'he3 : _GEN_1035; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1037 = 9'h1e4 == _T_215 ? 8'he4 : _GEN_1036; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1038 = 9'h1e5 == _T_215 ? 8'he5 : _GEN_1037; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1039 = 9'h1e6 == _T_215 ? 8'he6 : _GEN_1038; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1040 = 9'h1e7 == _T_215 ? 8'he7 : _GEN_1039; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1041 = 9'h1e8 == _T_215 ? 8'he8 : _GEN_1040; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1042 = 9'h1e9 == _T_215 ? 8'he9 : _GEN_1041; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1043 = 9'h1ea == _T_215 ? 8'hea : _GEN_1042; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1044 = 9'h1eb == _T_215 ? 8'heb : _GEN_1043; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1045 = 9'h1ec == _T_215 ? 8'hec : _GEN_1044; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1046 = 9'h1ed == _T_215 ? 8'hed : _GEN_1045; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1047 = 9'h1ee == _T_215 ? 8'hee : _GEN_1046; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1048 = 9'h1ef == _T_215 ? 8'hef : _GEN_1047; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1049 = 9'h1f0 == _T_215 ? 8'hf0 : _GEN_1048; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1050 = 9'h1f1 == _T_215 ? 8'hf1 : _GEN_1049; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1051 = 9'h1f2 == _T_215 ? 8'hf2 : _GEN_1050; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1052 = 9'h1f3 == _T_215 ? 8'hf3 : _GEN_1051; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1053 = 9'h1f4 == _T_215 ? 8'hf4 : _GEN_1052; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1054 = 9'h1f5 == _T_215 ? 8'hf5 : _GEN_1053; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1055 = 9'h1f6 == _T_215 ? 8'hf6 : _GEN_1054; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1056 = 9'h1f7 == _T_215 ? 8'hf7 : _GEN_1055; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1057 = 9'h1f8 == _T_215 ? 8'hf8 : _GEN_1056; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1058 = 9'h1f9 == _T_215 ? 8'hf9 : _GEN_1057; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1059 = 9'h1fa == _T_215 ? 8'hfa : _GEN_1058; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1060 = 9'h1fb == _T_215 ? 8'hfb : _GEN_1059; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1061 = 9'h1fc == _T_215 ? 8'hfc : _GEN_1060; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1062 = 9'h1fd == _T_215 ? 8'hfd : _GEN_1061; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1063 = 9'h1fe == _T_215 ? 8'hfe : _GEN_1062; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1064 = 9'h1ff == _T_215 ? 8'hff : _GEN_1063; // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1067 = 8'h1 == _GEN_1064 ? $signed(16'sh3fff) : $signed(16'sh4000); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1068 = 8'h1 == _GEN_1064 ? $signed(-16'shc9) : $signed(16'sh0); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1069 = 8'h2 == _GEN_1064 ? $signed(16'sh3ffb) : $signed(_GEN_1067); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1070 = 8'h2 == _GEN_1064 ? $signed(-16'sh192) : $signed(_GEN_1068); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1071 = 8'h3 == _GEN_1064 ? $signed(16'sh3ff5) : $signed(_GEN_1069); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1072 = 8'h3 == _GEN_1064 ? $signed(-16'sh25b) : $signed(_GEN_1070); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1073 = 8'h4 == _GEN_1064 ? $signed(16'sh3fec) : $signed(_GEN_1071); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1074 = 8'h4 == _GEN_1064 ? $signed(-16'sh324) : $signed(_GEN_1072); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1075 = 8'h5 == _GEN_1064 ? $signed(16'sh3fe1) : $signed(_GEN_1073); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1076 = 8'h5 == _GEN_1064 ? $signed(-16'sh3ed) : $signed(_GEN_1074); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1077 = 8'h6 == _GEN_1064 ? $signed(16'sh3fd4) : $signed(_GEN_1075); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1078 = 8'h6 == _GEN_1064 ? $signed(-16'sh4b5) : $signed(_GEN_1076); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1079 = 8'h7 == _GEN_1064 ? $signed(16'sh3fc4) : $signed(_GEN_1077); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1080 = 8'h7 == _GEN_1064 ? $signed(-16'sh57e) : $signed(_GEN_1078); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1081 = 8'h8 == _GEN_1064 ? $signed(16'sh3fb1) : $signed(_GEN_1079); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1082 = 8'h8 == _GEN_1064 ? $signed(-16'sh646) : $signed(_GEN_1080); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1083 = 8'h9 == _GEN_1064 ? $signed(16'sh3f9c) : $signed(_GEN_1081); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1084 = 8'h9 == _GEN_1064 ? $signed(-16'sh70e) : $signed(_GEN_1082); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1085 = 8'ha == _GEN_1064 ? $signed(16'sh3f85) : $signed(_GEN_1083); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1086 = 8'ha == _GEN_1064 ? $signed(-16'sh7d6) : $signed(_GEN_1084); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1087 = 8'hb == _GEN_1064 ? $signed(16'sh3f6b) : $signed(_GEN_1085); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1088 = 8'hb == _GEN_1064 ? $signed(-16'sh89d) : $signed(_GEN_1086); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1089 = 8'hc == _GEN_1064 ? $signed(16'sh3f4f) : $signed(_GEN_1087); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1090 = 8'hc == _GEN_1064 ? $signed(-16'sh964) : $signed(_GEN_1088); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1091 = 8'hd == _GEN_1064 ? $signed(16'sh3f30) : $signed(_GEN_1089); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1092 = 8'hd == _GEN_1064 ? $signed(-16'sha2b) : $signed(_GEN_1090); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1093 = 8'he == _GEN_1064 ? $signed(16'sh3f0f) : $signed(_GEN_1091); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1094 = 8'he == _GEN_1064 ? $signed(-16'shaf1) : $signed(_GEN_1092); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1095 = 8'hf == _GEN_1064 ? $signed(16'sh3eeb) : $signed(_GEN_1093); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1096 = 8'hf == _GEN_1064 ? $signed(-16'shbb7) : $signed(_GEN_1094); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1097 = 8'h10 == _GEN_1064 ? $signed(16'sh3ec5) : $signed(_GEN_1095); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1098 = 8'h10 == _GEN_1064 ? $signed(-16'shc7c) : $signed(_GEN_1096); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1099 = 8'h11 == _GEN_1064 ? $signed(16'sh3e9d) : $signed(_GEN_1097); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1100 = 8'h11 == _GEN_1064 ? $signed(-16'shd41) : $signed(_GEN_1098); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1101 = 8'h12 == _GEN_1064 ? $signed(16'sh3e72) : $signed(_GEN_1099); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1102 = 8'h12 == _GEN_1064 ? $signed(-16'she06) : $signed(_GEN_1100); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1103 = 8'h13 == _GEN_1064 ? $signed(16'sh3e45) : $signed(_GEN_1101); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1104 = 8'h13 == _GEN_1064 ? $signed(-16'sheca) : $signed(_GEN_1102); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1105 = 8'h14 == _GEN_1064 ? $signed(16'sh3e15) : $signed(_GEN_1103); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1106 = 8'h14 == _GEN_1064 ? $signed(-16'shf8d) : $signed(_GEN_1104); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1107 = 8'h15 == _GEN_1064 ? $signed(16'sh3de3) : $signed(_GEN_1105); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1108 = 8'h15 == _GEN_1064 ? $signed(-16'sh1050) : $signed(_GEN_1106); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1109 = 8'h16 == _GEN_1064 ? $signed(16'sh3daf) : $signed(_GEN_1107); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1110 = 8'h16 == _GEN_1064 ? $signed(-16'sh1112) : $signed(_GEN_1108); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1111 = 8'h17 == _GEN_1064 ? $signed(16'sh3d78) : $signed(_GEN_1109); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1112 = 8'h17 == _GEN_1064 ? $signed(-16'sh11d3) : $signed(_GEN_1110); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1113 = 8'h18 == _GEN_1064 ? $signed(16'sh3d3f) : $signed(_GEN_1111); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1114 = 8'h18 == _GEN_1064 ? $signed(-16'sh1294) : $signed(_GEN_1112); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1115 = 8'h19 == _GEN_1064 ? $signed(16'sh3d03) : $signed(_GEN_1113); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1116 = 8'h19 == _GEN_1064 ? $signed(-16'sh1354) : $signed(_GEN_1114); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1117 = 8'h1a == _GEN_1064 ? $signed(16'sh3cc5) : $signed(_GEN_1115); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1118 = 8'h1a == _GEN_1064 ? $signed(-16'sh1413) : $signed(_GEN_1116); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1119 = 8'h1b == _GEN_1064 ? $signed(16'sh3c85) : $signed(_GEN_1117); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1120 = 8'h1b == _GEN_1064 ? $signed(-16'sh14d2) : $signed(_GEN_1118); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1121 = 8'h1c == _GEN_1064 ? $signed(16'sh3c42) : $signed(_GEN_1119); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1122 = 8'h1c == _GEN_1064 ? $signed(-16'sh1590) : $signed(_GEN_1120); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1123 = 8'h1d == _GEN_1064 ? $signed(16'sh3bfd) : $signed(_GEN_1121); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1124 = 8'h1d == _GEN_1064 ? $signed(-16'sh164c) : $signed(_GEN_1122); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1125 = 8'h1e == _GEN_1064 ? $signed(16'sh3bb6) : $signed(_GEN_1123); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1126 = 8'h1e == _GEN_1064 ? $signed(-16'sh1709) : $signed(_GEN_1124); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1127 = 8'h1f == _GEN_1064 ? $signed(16'sh3b6d) : $signed(_GEN_1125); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1128 = 8'h1f == _GEN_1064 ? $signed(-16'sh17c4) : $signed(_GEN_1126); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1129 = 8'h20 == _GEN_1064 ? $signed(16'sh3b21) : $signed(_GEN_1127); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1130 = 8'h20 == _GEN_1064 ? $signed(-16'sh187e) : $signed(_GEN_1128); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1131 = 8'h21 == _GEN_1064 ? $signed(16'sh3ad3) : $signed(_GEN_1129); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1132 = 8'h21 == _GEN_1064 ? $signed(-16'sh1937) : $signed(_GEN_1130); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1133 = 8'h22 == _GEN_1064 ? $signed(16'sh3a82) : $signed(_GEN_1131); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1134 = 8'h22 == _GEN_1064 ? $signed(-16'sh19ef) : $signed(_GEN_1132); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1135 = 8'h23 == _GEN_1064 ? $signed(16'sh3a30) : $signed(_GEN_1133); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1136 = 8'h23 == _GEN_1064 ? $signed(-16'sh1aa7) : $signed(_GEN_1134); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1137 = 8'h24 == _GEN_1064 ? $signed(16'sh39db) : $signed(_GEN_1135); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1138 = 8'h24 == _GEN_1064 ? $signed(-16'sh1b5d) : $signed(_GEN_1136); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1139 = 8'h25 == _GEN_1064 ? $signed(16'sh3984) : $signed(_GEN_1137); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1140 = 8'h25 == _GEN_1064 ? $signed(-16'sh1c12) : $signed(_GEN_1138); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1141 = 8'h26 == _GEN_1064 ? $signed(16'sh392b) : $signed(_GEN_1139); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1142 = 8'h26 == _GEN_1064 ? $signed(-16'sh1cc6) : $signed(_GEN_1140); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1143 = 8'h27 == _GEN_1064 ? $signed(16'sh38cf) : $signed(_GEN_1141); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1144 = 8'h27 == _GEN_1064 ? $signed(-16'sh1d79) : $signed(_GEN_1142); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1145 = 8'h28 == _GEN_1064 ? $signed(16'sh3871) : $signed(_GEN_1143); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1146 = 8'h28 == _GEN_1064 ? $signed(-16'sh1e2b) : $signed(_GEN_1144); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1147 = 8'h29 == _GEN_1064 ? $signed(16'sh3812) : $signed(_GEN_1145); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1148 = 8'h29 == _GEN_1064 ? $signed(-16'sh1edc) : $signed(_GEN_1146); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1149 = 8'h2a == _GEN_1064 ? $signed(16'sh37b0) : $signed(_GEN_1147); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1150 = 8'h2a == _GEN_1064 ? $signed(-16'sh1f8c) : $signed(_GEN_1148); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1151 = 8'h2b == _GEN_1064 ? $signed(16'sh374b) : $signed(_GEN_1149); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1152 = 8'h2b == _GEN_1064 ? $signed(-16'sh203a) : $signed(_GEN_1150); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1153 = 8'h2c == _GEN_1064 ? $signed(16'sh36e5) : $signed(_GEN_1151); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1154 = 8'h2c == _GEN_1064 ? $signed(-16'sh20e7) : $signed(_GEN_1152); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1155 = 8'h2d == _GEN_1064 ? $signed(16'sh367d) : $signed(_GEN_1153); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1156 = 8'h2d == _GEN_1064 ? $signed(-16'sh2193) : $signed(_GEN_1154); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1157 = 8'h2e == _GEN_1064 ? $signed(16'sh3612) : $signed(_GEN_1155); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1158 = 8'h2e == _GEN_1064 ? $signed(-16'sh223d) : $signed(_GEN_1156); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1159 = 8'h2f == _GEN_1064 ? $signed(16'sh35a5) : $signed(_GEN_1157); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1160 = 8'h2f == _GEN_1064 ? $signed(-16'sh22e7) : $signed(_GEN_1158); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1161 = 8'h30 == _GEN_1064 ? $signed(16'sh3537) : $signed(_GEN_1159); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1162 = 8'h30 == _GEN_1064 ? $signed(-16'sh238e) : $signed(_GEN_1160); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1163 = 8'h31 == _GEN_1064 ? $signed(16'sh34c6) : $signed(_GEN_1161); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1164 = 8'h31 == _GEN_1064 ? $signed(-16'sh2435) : $signed(_GEN_1162); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1165 = 8'h32 == _GEN_1064 ? $signed(16'sh3453) : $signed(_GEN_1163); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1166 = 8'h32 == _GEN_1064 ? $signed(-16'sh24da) : $signed(_GEN_1164); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1167 = 8'h33 == _GEN_1064 ? $signed(16'sh33df) : $signed(_GEN_1165); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1168 = 8'h33 == _GEN_1064 ? $signed(-16'sh257e) : $signed(_GEN_1166); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1169 = 8'h34 == _GEN_1064 ? $signed(16'sh3368) : $signed(_GEN_1167); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1170 = 8'h34 == _GEN_1064 ? $signed(-16'sh2620) : $signed(_GEN_1168); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1171 = 8'h35 == _GEN_1064 ? $signed(16'sh32ef) : $signed(_GEN_1169); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1172 = 8'h35 == _GEN_1064 ? $signed(-16'sh26c1) : $signed(_GEN_1170); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1173 = 8'h36 == _GEN_1064 ? $signed(16'sh3274) : $signed(_GEN_1171); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1174 = 8'h36 == _GEN_1064 ? $signed(-16'sh2760) : $signed(_GEN_1172); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1175 = 8'h37 == _GEN_1064 ? $signed(16'sh31f8) : $signed(_GEN_1173); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1176 = 8'h37 == _GEN_1064 ? $signed(-16'sh27fe) : $signed(_GEN_1174); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1177 = 8'h38 == _GEN_1064 ? $signed(16'sh3179) : $signed(_GEN_1175); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1178 = 8'h38 == _GEN_1064 ? $signed(-16'sh289a) : $signed(_GEN_1176); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1179 = 8'h39 == _GEN_1064 ? $signed(16'sh30f9) : $signed(_GEN_1177); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1180 = 8'h39 == _GEN_1064 ? $signed(-16'sh2935) : $signed(_GEN_1178); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1181 = 8'h3a == _GEN_1064 ? $signed(16'sh3076) : $signed(_GEN_1179); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1182 = 8'h3a == _GEN_1064 ? $signed(-16'sh29ce) : $signed(_GEN_1180); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1183 = 8'h3b == _GEN_1064 ? $signed(16'sh2ff2) : $signed(_GEN_1181); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1184 = 8'h3b == _GEN_1064 ? $signed(-16'sh2a65) : $signed(_GEN_1182); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1185 = 8'h3c == _GEN_1064 ? $signed(16'sh2f6c) : $signed(_GEN_1183); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1186 = 8'h3c == _GEN_1064 ? $signed(-16'sh2afb) : $signed(_GEN_1184); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1187 = 8'h3d == _GEN_1064 ? $signed(16'sh2ee4) : $signed(_GEN_1185); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1188 = 8'h3d == _GEN_1064 ? $signed(-16'sh2b8f) : $signed(_GEN_1186); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1189 = 8'h3e == _GEN_1064 ? $signed(16'sh2e5a) : $signed(_GEN_1187); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1190 = 8'h3e == _GEN_1064 ? $signed(-16'sh2c21) : $signed(_GEN_1188); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1191 = 8'h3f == _GEN_1064 ? $signed(16'sh2dcf) : $signed(_GEN_1189); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1192 = 8'h3f == _GEN_1064 ? $signed(-16'sh2cb2) : $signed(_GEN_1190); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1193 = 8'h40 == _GEN_1064 ? $signed(16'sh2d41) : $signed(_GEN_1191); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1194 = 8'h40 == _GEN_1064 ? $signed(-16'sh2d41) : $signed(_GEN_1192); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1195 = 8'h41 == _GEN_1064 ? $signed(16'sh2cb2) : $signed(_GEN_1193); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1196 = 8'h41 == _GEN_1064 ? $signed(-16'sh2dcf) : $signed(_GEN_1194); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1197 = 8'h42 == _GEN_1064 ? $signed(16'sh2c21) : $signed(_GEN_1195); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1198 = 8'h42 == _GEN_1064 ? $signed(-16'sh2e5a) : $signed(_GEN_1196); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1199 = 8'h43 == _GEN_1064 ? $signed(16'sh2b8f) : $signed(_GEN_1197); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1200 = 8'h43 == _GEN_1064 ? $signed(-16'sh2ee4) : $signed(_GEN_1198); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1201 = 8'h44 == _GEN_1064 ? $signed(16'sh2afb) : $signed(_GEN_1199); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1202 = 8'h44 == _GEN_1064 ? $signed(-16'sh2f6c) : $signed(_GEN_1200); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1203 = 8'h45 == _GEN_1064 ? $signed(16'sh2a65) : $signed(_GEN_1201); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1204 = 8'h45 == _GEN_1064 ? $signed(-16'sh2ff2) : $signed(_GEN_1202); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1205 = 8'h46 == _GEN_1064 ? $signed(16'sh29ce) : $signed(_GEN_1203); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1206 = 8'h46 == _GEN_1064 ? $signed(-16'sh3076) : $signed(_GEN_1204); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1207 = 8'h47 == _GEN_1064 ? $signed(16'sh2935) : $signed(_GEN_1205); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1208 = 8'h47 == _GEN_1064 ? $signed(-16'sh30f9) : $signed(_GEN_1206); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1209 = 8'h48 == _GEN_1064 ? $signed(16'sh289a) : $signed(_GEN_1207); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1210 = 8'h48 == _GEN_1064 ? $signed(-16'sh3179) : $signed(_GEN_1208); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1211 = 8'h49 == _GEN_1064 ? $signed(16'sh27fe) : $signed(_GEN_1209); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1212 = 8'h49 == _GEN_1064 ? $signed(-16'sh31f8) : $signed(_GEN_1210); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1213 = 8'h4a == _GEN_1064 ? $signed(16'sh2760) : $signed(_GEN_1211); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1214 = 8'h4a == _GEN_1064 ? $signed(-16'sh3274) : $signed(_GEN_1212); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1215 = 8'h4b == _GEN_1064 ? $signed(16'sh26c1) : $signed(_GEN_1213); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1216 = 8'h4b == _GEN_1064 ? $signed(-16'sh32ef) : $signed(_GEN_1214); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1217 = 8'h4c == _GEN_1064 ? $signed(16'sh2620) : $signed(_GEN_1215); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1218 = 8'h4c == _GEN_1064 ? $signed(-16'sh3368) : $signed(_GEN_1216); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1219 = 8'h4d == _GEN_1064 ? $signed(16'sh257e) : $signed(_GEN_1217); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1220 = 8'h4d == _GEN_1064 ? $signed(-16'sh33df) : $signed(_GEN_1218); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1221 = 8'h4e == _GEN_1064 ? $signed(16'sh24da) : $signed(_GEN_1219); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1222 = 8'h4e == _GEN_1064 ? $signed(-16'sh3453) : $signed(_GEN_1220); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1223 = 8'h4f == _GEN_1064 ? $signed(16'sh2435) : $signed(_GEN_1221); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1224 = 8'h4f == _GEN_1064 ? $signed(-16'sh34c6) : $signed(_GEN_1222); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1225 = 8'h50 == _GEN_1064 ? $signed(16'sh238e) : $signed(_GEN_1223); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1226 = 8'h50 == _GEN_1064 ? $signed(-16'sh3537) : $signed(_GEN_1224); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1227 = 8'h51 == _GEN_1064 ? $signed(16'sh22e7) : $signed(_GEN_1225); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1228 = 8'h51 == _GEN_1064 ? $signed(-16'sh35a5) : $signed(_GEN_1226); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1229 = 8'h52 == _GEN_1064 ? $signed(16'sh223d) : $signed(_GEN_1227); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1230 = 8'h52 == _GEN_1064 ? $signed(-16'sh3612) : $signed(_GEN_1228); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1231 = 8'h53 == _GEN_1064 ? $signed(16'sh2193) : $signed(_GEN_1229); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1232 = 8'h53 == _GEN_1064 ? $signed(-16'sh367d) : $signed(_GEN_1230); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1233 = 8'h54 == _GEN_1064 ? $signed(16'sh20e7) : $signed(_GEN_1231); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1234 = 8'h54 == _GEN_1064 ? $signed(-16'sh36e5) : $signed(_GEN_1232); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1235 = 8'h55 == _GEN_1064 ? $signed(16'sh203a) : $signed(_GEN_1233); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1236 = 8'h55 == _GEN_1064 ? $signed(-16'sh374b) : $signed(_GEN_1234); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1237 = 8'h56 == _GEN_1064 ? $signed(16'sh1f8c) : $signed(_GEN_1235); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1238 = 8'h56 == _GEN_1064 ? $signed(-16'sh37b0) : $signed(_GEN_1236); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1239 = 8'h57 == _GEN_1064 ? $signed(16'sh1edc) : $signed(_GEN_1237); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1240 = 8'h57 == _GEN_1064 ? $signed(-16'sh3812) : $signed(_GEN_1238); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1241 = 8'h58 == _GEN_1064 ? $signed(16'sh1e2b) : $signed(_GEN_1239); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1242 = 8'h58 == _GEN_1064 ? $signed(-16'sh3871) : $signed(_GEN_1240); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1243 = 8'h59 == _GEN_1064 ? $signed(16'sh1d79) : $signed(_GEN_1241); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1244 = 8'h59 == _GEN_1064 ? $signed(-16'sh38cf) : $signed(_GEN_1242); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1245 = 8'h5a == _GEN_1064 ? $signed(16'sh1cc6) : $signed(_GEN_1243); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1246 = 8'h5a == _GEN_1064 ? $signed(-16'sh392b) : $signed(_GEN_1244); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1247 = 8'h5b == _GEN_1064 ? $signed(16'sh1c12) : $signed(_GEN_1245); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1248 = 8'h5b == _GEN_1064 ? $signed(-16'sh3984) : $signed(_GEN_1246); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1249 = 8'h5c == _GEN_1064 ? $signed(16'sh1b5d) : $signed(_GEN_1247); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1250 = 8'h5c == _GEN_1064 ? $signed(-16'sh39db) : $signed(_GEN_1248); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1251 = 8'h5d == _GEN_1064 ? $signed(16'sh1aa7) : $signed(_GEN_1249); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1252 = 8'h5d == _GEN_1064 ? $signed(-16'sh3a30) : $signed(_GEN_1250); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1253 = 8'h5e == _GEN_1064 ? $signed(16'sh19ef) : $signed(_GEN_1251); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1254 = 8'h5e == _GEN_1064 ? $signed(-16'sh3a82) : $signed(_GEN_1252); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1255 = 8'h5f == _GEN_1064 ? $signed(16'sh1937) : $signed(_GEN_1253); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1256 = 8'h5f == _GEN_1064 ? $signed(-16'sh3ad3) : $signed(_GEN_1254); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1257 = 8'h60 == _GEN_1064 ? $signed(16'sh187e) : $signed(_GEN_1255); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1258 = 8'h60 == _GEN_1064 ? $signed(-16'sh3b21) : $signed(_GEN_1256); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1259 = 8'h61 == _GEN_1064 ? $signed(16'sh17c4) : $signed(_GEN_1257); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1260 = 8'h61 == _GEN_1064 ? $signed(-16'sh3b6d) : $signed(_GEN_1258); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1261 = 8'h62 == _GEN_1064 ? $signed(16'sh1709) : $signed(_GEN_1259); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1262 = 8'h62 == _GEN_1064 ? $signed(-16'sh3bb6) : $signed(_GEN_1260); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1263 = 8'h63 == _GEN_1064 ? $signed(16'sh164c) : $signed(_GEN_1261); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1264 = 8'h63 == _GEN_1064 ? $signed(-16'sh3bfd) : $signed(_GEN_1262); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1265 = 8'h64 == _GEN_1064 ? $signed(16'sh1590) : $signed(_GEN_1263); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1266 = 8'h64 == _GEN_1064 ? $signed(-16'sh3c42) : $signed(_GEN_1264); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1267 = 8'h65 == _GEN_1064 ? $signed(16'sh14d2) : $signed(_GEN_1265); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1268 = 8'h65 == _GEN_1064 ? $signed(-16'sh3c85) : $signed(_GEN_1266); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1269 = 8'h66 == _GEN_1064 ? $signed(16'sh1413) : $signed(_GEN_1267); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1270 = 8'h66 == _GEN_1064 ? $signed(-16'sh3cc5) : $signed(_GEN_1268); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1271 = 8'h67 == _GEN_1064 ? $signed(16'sh1354) : $signed(_GEN_1269); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1272 = 8'h67 == _GEN_1064 ? $signed(-16'sh3d03) : $signed(_GEN_1270); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1273 = 8'h68 == _GEN_1064 ? $signed(16'sh1294) : $signed(_GEN_1271); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1274 = 8'h68 == _GEN_1064 ? $signed(-16'sh3d3f) : $signed(_GEN_1272); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1275 = 8'h69 == _GEN_1064 ? $signed(16'sh11d3) : $signed(_GEN_1273); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1276 = 8'h69 == _GEN_1064 ? $signed(-16'sh3d78) : $signed(_GEN_1274); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1277 = 8'h6a == _GEN_1064 ? $signed(16'sh1112) : $signed(_GEN_1275); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1278 = 8'h6a == _GEN_1064 ? $signed(-16'sh3daf) : $signed(_GEN_1276); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1279 = 8'h6b == _GEN_1064 ? $signed(16'sh1050) : $signed(_GEN_1277); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1280 = 8'h6b == _GEN_1064 ? $signed(-16'sh3de3) : $signed(_GEN_1278); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1281 = 8'h6c == _GEN_1064 ? $signed(16'shf8d) : $signed(_GEN_1279); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1282 = 8'h6c == _GEN_1064 ? $signed(-16'sh3e15) : $signed(_GEN_1280); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1283 = 8'h6d == _GEN_1064 ? $signed(16'sheca) : $signed(_GEN_1281); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1284 = 8'h6d == _GEN_1064 ? $signed(-16'sh3e45) : $signed(_GEN_1282); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1285 = 8'h6e == _GEN_1064 ? $signed(16'she06) : $signed(_GEN_1283); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1286 = 8'h6e == _GEN_1064 ? $signed(-16'sh3e72) : $signed(_GEN_1284); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1287 = 8'h6f == _GEN_1064 ? $signed(16'shd41) : $signed(_GEN_1285); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1288 = 8'h6f == _GEN_1064 ? $signed(-16'sh3e9d) : $signed(_GEN_1286); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1289 = 8'h70 == _GEN_1064 ? $signed(16'shc7c) : $signed(_GEN_1287); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1290 = 8'h70 == _GEN_1064 ? $signed(-16'sh3ec5) : $signed(_GEN_1288); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1291 = 8'h71 == _GEN_1064 ? $signed(16'shbb7) : $signed(_GEN_1289); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1292 = 8'h71 == _GEN_1064 ? $signed(-16'sh3eeb) : $signed(_GEN_1290); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1293 = 8'h72 == _GEN_1064 ? $signed(16'shaf1) : $signed(_GEN_1291); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1294 = 8'h72 == _GEN_1064 ? $signed(-16'sh3f0f) : $signed(_GEN_1292); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1295 = 8'h73 == _GEN_1064 ? $signed(16'sha2b) : $signed(_GEN_1293); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1296 = 8'h73 == _GEN_1064 ? $signed(-16'sh3f30) : $signed(_GEN_1294); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1297 = 8'h74 == _GEN_1064 ? $signed(16'sh964) : $signed(_GEN_1295); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1298 = 8'h74 == _GEN_1064 ? $signed(-16'sh3f4f) : $signed(_GEN_1296); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1299 = 8'h75 == _GEN_1064 ? $signed(16'sh89d) : $signed(_GEN_1297); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1300 = 8'h75 == _GEN_1064 ? $signed(-16'sh3f6b) : $signed(_GEN_1298); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1301 = 8'h76 == _GEN_1064 ? $signed(16'sh7d6) : $signed(_GEN_1299); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1302 = 8'h76 == _GEN_1064 ? $signed(-16'sh3f85) : $signed(_GEN_1300); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1303 = 8'h77 == _GEN_1064 ? $signed(16'sh70e) : $signed(_GEN_1301); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1304 = 8'h77 == _GEN_1064 ? $signed(-16'sh3f9c) : $signed(_GEN_1302); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1305 = 8'h78 == _GEN_1064 ? $signed(16'sh646) : $signed(_GEN_1303); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1306 = 8'h78 == _GEN_1064 ? $signed(-16'sh3fb1) : $signed(_GEN_1304); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1307 = 8'h79 == _GEN_1064 ? $signed(16'sh57e) : $signed(_GEN_1305); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1308 = 8'h79 == _GEN_1064 ? $signed(-16'sh3fc4) : $signed(_GEN_1306); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1309 = 8'h7a == _GEN_1064 ? $signed(16'sh4b5) : $signed(_GEN_1307); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1310 = 8'h7a == _GEN_1064 ? $signed(-16'sh3fd4) : $signed(_GEN_1308); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1311 = 8'h7b == _GEN_1064 ? $signed(16'sh3ed) : $signed(_GEN_1309); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1312 = 8'h7b == _GEN_1064 ? $signed(-16'sh3fe1) : $signed(_GEN_1310); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1313 = 8'h7c == _GEN_1064 ? $signed(16'sh324) : $signed(_GEN_1311); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1314 = 8'h7c == _GEN_1064 ? $signed(-16'sh3fec) : $signed(_GEN_1312); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1315 = 8'h7d == _GEN_1064 ? $signed(16'sh25b) : $signed(_GEN_1313); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1316 = 8'h7d == _GEN_1064 ? $signed(-16'sh3ff5) : $signed(_GEN_1314); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1317 = 8'h7e == _GEN_1064 ? $signed(16'sh192) : $signed(_GEN_1315); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1318 = 8'h7e == _GEN_1064 ? $signed(-16'sh3ffb) : $signed(_GEN_1316); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1319 = 8'h7f == _GEN_1064 ? $signed(16'shc9) : $signed(_GEN_1317); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1320 = 8'h7f == _GEN_1064 ? $signed(-16'sh3fff) : $signed(_GEN_1318); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1321 = 8'h80 == _GEN_1064 ? $signed(16'sh0) : $signed(_GEN_1319); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1322 = 8'h80 == _GEN_1064 ? $signed(-16'sh4000) : $signed(_GEN_1320); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1323 = 8'h81 == _GEN_1064 ? $signed(-16'shc9) : $signed(_GEN_1321); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1324 = 8'h81 == _GEN_1064 ? $signed(-16'sh3fff) : $signed(_GEN_1322); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1325 = 8'h82 == _GEN_1064 ? $signed(-16'sh192) : $signed(_GEN_1323); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1326 = 8'h82 == _GEN_1064 ? $signed(-16'sh3ffb) : $signed(_GEN_1324); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1327 = 8'h83 == _GEN_1064 ? $signed(-16'sh324) : $signed(_GEN_1325); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1328 = 8'h83 == _GEN_1064 ? $signed(-16'sh3fec) : $signed(_GEN_1326); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1329 = 8'h84 == _GEN_1064 ? $signed(-16'sh4b5) : $signed(_GEN_1327); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1330 = 8'h84 == _GEN_1064 ? $signed(-16'sh3fd4) : $signed(_GEN_1328); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1331 = 8'h85 == _GEN_1064 ? $signed(-16'sh57e) : $signed(_GEN_1329); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1332 = 8'h85 == _GEN_1064 ? $signed(-16'sh3fc4) : $signed(_GEN_1330); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1333 = 8'h86 == _GEN_1064 ? $signed(-16'sh646) : $signed(_GEN_1331); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1334 = 8'h86 == _GEN_1064 ? $signed(-16'sh3fb1) : $signed(_GEN_1332); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1335 = 8'h87 == _GEN_1064 ? $signed(-16'sh7d6) : $signed(_GEN_1333); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1336 = 8'h87 == _GEN_1064 ? $signed(-16'sh3f85) : $signed(_GEN_1334); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1337 = 8'h88 == _GEN_1064 ? $signed(-16'sh964) : $signed(_GEN_1335); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1338 = 8'h88 == _GEN_1064 ? $signed(-16'sh3f4f) : $signed(_GEN_1336); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1339 = 8'h89 == _GEN_1064 ? $signed(-16'sha2b) : $signed(_GEN_1337); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1340 = 8'h89 == _GEN_1064 ? $signed(-16'sh3f30) : $signed(_GEN_1338); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1341 = 8'h8a == _GEN_1064 ? $signed(-16'shaf1) : $signed(_GEN_1339); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1342 = 8'h8a == _GEN_1064 ? $signed(-16'sh3f0f) : $signed(_GEN_1340); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1343 = 8'h8b == _GEN_1064 ? $signed(-16'shc7c) : $signed(_GEN_1341); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1344 = 8'h8b == _GEN_1064 ? $signed(-16'sh3ec5) : $signed(_GEN_1342); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1345 = 8'h8c == _GEN_1064 ? $signed(-16'she06) : $signed(_GEN_1343); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1346 = 8'h8c == _GEN_1064 ? $signed(-16'sh3e72) : $signed(_GEN_1344); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1347 = 8'h8d == _GEN_1064 ? $signed(-16'sheca) : $signed(_GEN_1345); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1348 = 8'h8d == _GEN_1064 ? $signed(-16'sh3e45) : $signed(_GEN_1346); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1349 = 8'h8e == _GEN_1064 ? $signed(-16'shf8d) : $signed(_GEN_1347); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1350 = 8'h8e == _GEN_1064 ? $signed(-16'sh3e15) : $signed(_GEN_1348); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1351 = 8'h8f == _GEN_1064 ? $signed(-16'sh1112) : $signed(_GEN_1349); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1352 = 8'h8f == _GEN_1064 ? $signed(-16'sh3daf) : $signed(_GEN_1350); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1353 = 8'h90 == _GEN_1064 ? $signed(-16'sh1294) : $signed(_GEN_1351); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1354 = 8'h90 == _GEN_1064 ? $signed(-16'sh3d3f) : $signed(_GEN_1352); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1355 = 8'h91 == _GEN_1064 ? $signed(-16'sh1354) : $signed(_GEN_1353); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1356 = 8'h91 == _GEN_1064 ? $signed(-16'sh3d03) : $signed(_GEN_1354); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1357 = 8'h92 == _GEN_1064 ? $signed(-16'sh1413) : $signed(_GEN_1355); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1358 = 8'h92 == _GEN_1064 ? $signed(-16'sh3cc5) : $signed(_GEN_1356); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1359 = 8'h93 == _GEN_1064 ? $signed(-16'sh1590) : $signed(_GEN_1357); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1360 = 8'h93 == _GEN_1064 ? $signed(-16'sh3c42) : $signed(_GEN_1358); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1361 = 8'h94 == _GEN_1064 ? $signed(-16'sh1709) : $signed(_GEN_1359); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1362 = 8'h94 == _GEN_1064 ? $signed(-16'sh3bb6) : $signed(_GEN_1360); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1363 = 8'h95 == _GEN_1064 ? $signed(-16'sh17c4) : $signed(_GEN_1361); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1364 = 8'h95 == _GEN_1064 ? $signed(-16'sh3b6d) : $signed(_GEN_1362); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1365 = 8'h96 == _GEN_1064 ? $signed(-16'sh187e) : $signed(_GEN_1363); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1366 = 8'h96 == _GEN_1064 ? $signed(-16'sh3b21) : $signed(_GEN_1364); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1367 = 8'h97 == _GEN_1064 ? $signed(-16'sh19ef) : $signed(_GEN_1365); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1368 = 8'h97 == _GEN_1064 ? $signed(-16'sh3a82) : $signed(_GEN_1366); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1369 = 8'h98 == _GEN_1064 ? $signed(-16'sh1b5d) : $signed(_GEN_1367); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1370 = 8'h98 == _GEN_1064 ? $signed(-16'sh39db) : $signed(_GEN_1368); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1371 = 8'h99 == _GEN_1064 ? $signed(-16'sh1c12) : $signed(_GEN_1369); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1372 = 8'h99 == _GEN_1064 ? $signed(-16'sh3984) : $signed(_GEN_1370); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1373 = 8'h9a == _GEN_1064 ? $signed(-16'sh1cc6) : $signed(_GEN_1371); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1374 = 8'h9a == _GEN_1064 ? $signed(-16'sh392b) : $signed(_GEN_1372); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1375 = 8'h9b == _GEN_1064 ? $signed(-16'sh1e2b) : $signed(_GEN_1373); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1376 = 8'h9b == _GEN_1064 ? $signed(-16'sh3871) : $signed(_GEN_1374); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1377 = 8'h9c == _GEN_1064 ? $signed(-16'sh1f8c) : $signed(_GEN_1375); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1378 = 8'h9c == _GEN_1064 ? $signed(-16'sh37b0) : $signed(_GEN_1376); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1379 = 8'h9d == _GEN_1064 ? $signed(-16'sh203a) : $signed(_GEN_1377); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1380 = 8'h9d == _GEN_1064 ? $signed(-16'sh374b) : $signed(_GEN_1378); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1381 = 8'h9e == _GEN_1064 ? $signed(-16'sh20e7) : $signed(_GEN_1379); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1382 = 8'h9e == _GEN_1064 ? $signed(-16'sh36e5) : $signed(_GEN_1380); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1383 = 8'h9f == _GEN_1064 ? $signed(-16'sh223d) : $signed(_GEN_1381); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1384 = 8'h9f == _GEN_1064 ? $signed(-16'sh3612) : $signed(_GEN_1382); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1385 = 8'ha0 == _GEN_1064 ? $signed(-16'sh238e) : $signed(_GEN_1383); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1386 = 8'ha0 == _GEN_1064 ? $signed(-16'sh3537) : $signed(_GEN_1384); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1387 = 8'ha1 == _GEN_1064 ? $signed(-16'sh2435) : $signed(_GEN_1385); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1388 = 8'ha1 == _GEN_1064 ? $signed(-16'sh34c6) : $signed(_GEN_1386); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1389 = 8'ha2 == _GEN_1064 ? $signed(-16'sh24da) : $signed(_GEN_1387); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1390 = 8'ha2 == _GEN_1064 ? $signed(-16'sh3453) : $signed(_GEN_1388); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1391 = 8'ha3 == _GEN_1064 ? $signed(-16'sh2620) : $signed(_GEN_1389); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1392 = 8'ha3 == _GEN_1064 ? $signed(-16'sh3368) : $signed(_GEN_1390); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1393 = 8'ha4 == _GEN_1064 ? $signed(-16'sh2760) : $signed(_GEN_1391); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1394 = 8'ha4 == _GEN_1064 ? $signed(-16'sh3274) : $signed(_GEN_1392); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1395 = 8'ha5 == _GEN_1064 ? $signed(-16'sh27fe) : $signed(_GEN_1393); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1396 = 8'ha5 == _GEN_1064 ? $signed(-16'sh31f8) : $signed(_GEN_1394); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1397 = 8'ha6 == _GEN_1064 ? $signed(-16'sh289a) : $signed(_GEN_1395); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1398 = 8'ha6 == _GEN_1064 ? $signed(-16'sh3179) : $signed(_GEN_1396); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1399 = 8'ha7 == _GEN_1064 ? $signed(-16'sh29ce) : $signed(_GEN_1397); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1400 = 8'ha7 == _GEN_1064 ? $signed(-16'sh3076) : $signed(_GEN_1398); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1401 = 8'ha8 == _GEN_1064 ? $signed(-16'sh2afb) : $signed(_GEN_1399); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1402 = 8'ha8 == _GEN_1064 ? $signed(-16'sh2f6c) : $signed(_GEN_1400); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1403 = 8'ha9 == _GEN_1064 ? $signed(-16'sh2b8f) : $signed(_GEN_1401); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1404 = 8'ha9 == _GEN_1064 ? $signed(-16'sh2ee4) : $signed(_GEN_1402); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1405 = 8'haa == _GEN_1064 ? $signed(-16'sh2c21) : $signed(_GEN_1403); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1406 = 8'haa == _GEN_1064 ? $signed(-16'sh2e5a) : $signed(_GEN_1404); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1407 = 8'hab == _GEN_1064 ? $signed(-16'sh2d41) : $signed(_GEN_1405); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1408 = 8'hab == _GEN_1064 ? $signed(-16'sh2d41) : $signed(_GEN_1406); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1409 = 8'hac == _GEN_1064 ? $signed(-16'sh2e5a) : $signed(_GEN_1407); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1410 = 8'hac == _GEN_1064 ? $signed(-16'sh2c21) : $signed(_GEN_1408); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1411 = 8'had == _GEN_1064 ? $signed(-16'sh2ee4) : $signed(_GEN_1409); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1412 = 8'had == _GEN_1064 ? $signed(-16'sh2b8f) : $signed(_GEN_1410); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1413 = 8'hae == _GEN_1064 ? $signed(-16'sh2f6c) : $signed(_GEN_1411); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1414 = 8'hae == _GEN_1064 ? $signed(-16'sh2afb) : $signed(_GEN_1412); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1415 = 8'haf == _GEN_1064 ? $signed(-16'sh3076) : $signed(_GEN_1413); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1416 = 8'haf == _GEN_1064 ? $signed(-16'sh29ce) : $signed(_GEN_1414); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1417 = 8'hb0 == _GEN_1064 ? $signed(-16'sh3179) : $signed(_GEN_1415); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1418 = 8'hb0 == _GEN_1064 ? $signed(-16'sh289a) : $signed(_GEN_1416); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1419 = 8'hb1 == _GEN_1064 ? $signed(-16'sh31f8) : $signed(_GEN_1417); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1420 = 8'hb1 == _GEN_1064 ? $signed(-16'sh27fe) : $signed(_GEN_1418); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1421 = 8'hb2 == _GEN_1064 ? $signed(-16'sh3274) : $signed(_GEN_1419); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1422 = 8'hb2 == _GEN_1064 ? $signed(-16'sh2760) : $signed(_GEN_1420); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1423 = 8'hb3 == _GEN_1064 ? $signed(-16'sh3368) : $signed(_GEN_1421); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1424 = 8'hb3 == _GEN_1064 ? $signed(-16'sh2620) : $signed(_GEN_1422); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1425 = 8'hb4 == _GEN_1064 ? $signed(-16'sh3453) : $signed(_GEN_1423); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1426 = 8'hb4 == _GEN_1064 ? $signed(-16'sh24da) : $signed(_GEN_1424); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1427 = 8'hb5 == _GEN_1064 ? $signed(-16'sh34c6) : $signed(_GEN_1425); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1428 = 8'hb5 == _GEN_1064 ? $signed(-16'sh2435) : $signed(_GEN_1426); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1429 = 8'hb6 == _GEN_1064 ? $signed(-16'sh3537) : $signed(_GEN_1427); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1430 = 8'hb6 == _GEN_1064 ? $signed(-16'sh238e) : $signed(_GEN_1428); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1431 = 8'hb7 == _GEN_1064 ? $signed(-16'sh3612) : $signed(_GEN_1429); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1432 = 8'hb7 == _GEN_1064 ? $signed(-16'sh223d) : $signed(_GEN_1430); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1433 = 8'hb8 == _GEN_1064 ? $signed(-16'sh36e5) : $signed(_GEN_1431); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1434 = 8'hb8 == _GEN_1064 ? $signed(-16'sh20e7) : $signed(_GEN_1432); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1435 = 8'hb9 == _GEN_1064 ? $signed(-16'sh374b) : $signed(_GEN_1433); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1436 = 8'hb9 == _GEN_1064 ? $signed(-16'sh203a) : $signed(_GEN_1434); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1437 = 8'hba == _GEN_1064 ? $signed(-16'sh37b0) : $signed(_GEN_1435); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1438 = 8'hba == _GEN_1064 ? $signed(-16'sh1f8c) : $signed(_GEN_1436); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1439 = 8'hbb == _GEN_1064 ? $signed(-16'sh3871) : $signed(_GEN_1437); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1440 = 8'hbb == _GEN_1064 ? $signed(-16'sh1e2b) : $signed(_GEN_1438); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1441 = 8'hbc == _GEN_1064 ? $signed(-16'sh392b) : $signed(_GEN_1439); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1442 = 8'hbc == _GEN_1064 ? $signed(-16'sh1cc6) : $signed(_GEN_1440); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1443 = 8'hbd == _GEN_1064 ? $signed(-16'sh3984) : $signed(_GEN_1441); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1444 = 8'hbd == _GEN_1064 ? $signed(-16'sh1c12) : $signed(_GEN_1442); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1445 = 8'hbe == _GEN_1064 ? $signed(-16'sh39db) : $signed(_GEN_1443); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1446 = 8'hbe == _GEN_1064 ? $signed(-16'sh1b5d) : $signed(_GEN_1444); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1447 = 8'hbf == _GEN_1064 ? $signed(-16'sh3a82) : $signed(_GEN_1445); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1448 = 8'hbf == _GEN_1064 ? $signed(-16'sh19ef) : $signed(_GEN_1446); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1449 = 8'hc0 == _GEN_1064 ? $signed(-16'sh3b21) : $signed(_GEN_1447); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1450 = 8'hc0 == _GEN_1064 ? $signed(-16'sh187e) : $signed(_GEN_1448); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1451 = 8'hc1 == _GEN_1064 ? $signed(-16'sh3b6d) : $signed(_GEN_1449); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1452 = 8'hc1 == _GEN_1064 ? $signed(-16'sh17c4) : $signed(_GEN_1450); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1453 = 8'hc2 == _GEN_1064 ? $signed(-16'sh3bb6) : $signed(_GEN_1451); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1454 = 8'hc2 == _GEN_1064 ? $signed(-16'sh1709) : $signed(_GEN_1452); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1455 = 8'hc3 == _GEN_1064 ? $signed(-16'sh3c42) : $signed(_GEN_1453); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1456 = 8'hc3 == _GEN_1064 ? $signed(-16'sh1590) : $signed(_GEN_1454); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1457 = 8'hc4 == _GEN_1064 ? $signed(-16'sh3cc5) : $signed(_GEN_1455); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1458 = 8'hc4 == _GEN_1064 ? $signed(-16'sh1413) : $signed(_GEN_1456); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1459 = 8'hc5 == _GEN_1064 ? $signed(-16'sh3d03) : $signed(_GEN_1457); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1460 = 8'hc5 == _GEN_1064 ? $signed(-16'sh1354) : $signed(_GEN_1458); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1461 = 8'hc6 == _GEN_1064 ? $signed(-16'sh3d3f) : $signed(_GEN_1459); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1462 = 8'hc6 == _GEN_1064 ? $signed(-16'sh1294) : $signed(_GEN_1460); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1463 = 8'hc7 == _GEN_1064 ? $signed(-16'sh3daf) : $signed(_GEN_1461); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1464 = 8'hc7 == _GEN_1064 ? $signed(-16'sh1112) : $signed(_GEN_1462); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1465 = 8'hc8 == _GEN_1064 ? $signed(-16'sh3e15) : $signed(_GEN_1463); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1466 = 8'hc8 == _GEN_1064 ? $signed(-16'shf8d) : $signed(_GEN_1464); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1467 = 8'hc9 == _GEN_1064 ? $signed(-16'sh3e45) : $signed(_GEN_1465); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1468 = 8'hc9 == _GEN_1064 ? $signed(-16'sheca) : $signed(_GEN_1466); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1469 = 8'hca == _GEN_1064 ? $signed(-16'sh3e72) : $signed(_GEN_1467); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1470 = 8'hca == _GEN_1064 ? $signed(-16'she06) : $signed(_GEN_1468); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1471 = 8'hcb == _GEN_1064 ? $signed(-16'sh3ec5) : $signed(_GEN_1469); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1472 = 8'hcb == _GEN_1064 ? $signed(-16'shc7c) : $signed(_GEN_1470); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1473 = 8'hcc == _GEN_1064 ? $signed(-16'sh3f0f) : $signed(_GEN_1471); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1474 = 8'hcc == _GEN_1064 ? $signed(-16'shaf1) : $signed(_GEN_1472); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1475 = 8'hcd == _GEN_1064 ? $signed(-16'sh3f30) : $signed(_GEN_1473); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1476 = 8'hcd == _GEN_1064 ? $signed(-16'sha2b) : $signed(_GEN_1474); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1477 = 8'hce == _GEN_1064 ? $signed(-16'sh3f4f) : $signed(_GEN_1475); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1478 = 8'hce == _GEN_1064 ? $signed(-16'sh964) : $signed(_GEN_1476); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1479 = 8'hcf == _GEN_1064 ? $signed(-16'sh3f85) : $signed(_GEN_1477); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1480 = 8'hcf == _GEN_1064 ? $signed(-16'sh7d6) : $signed(_GEN_1478); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1481 = 8'hd0 == _GEN_1064 ? $signed(-16'sh3fb1) : $signed(_GEN_1479); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1482 = 8'hd0 == _GEN_1064 ? $signed(-16'sh646) : $signed(_GEN_1480); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1483 = 8'hd1 == _GEN_1064 ? $signed(-16'sh3fc4) : $signed(_GEN_1481); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1484 = 8'hd1 == _GEN_1064 ? $signed(-16'sh57e) : $signed(_GEN_1482); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1485 = 8'hd2 == _GEN_1064 ? $signed(-16'sh3fd4) : $signed(_GEN_1483); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1486 = 8'hd2 == _GEN_1064 ? $signed(-16'sh4b5) : $signed(_GEN_1484); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1487 = 8'hd3 == _GEN_1064 ? $signed(-16'sh3fec) : $signed(_GEN_1485); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1488 = 8'hd3 == _GEN_1064 ? $signed(-16'sh324) : $signed(_GEN_1486); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1489 = 8'hd4 == _GEN_1064 ? $signed(-16'sh3ffb) : $signed(_GEN_1487); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1490 = 8'hd4 == _GEN_1064 ? $signed(-16'sh192) : $signed(_GEN_1488); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1491 = 8'hd5 == _GEN_1064 ? $signed(-16'sh3fff) : $signed(_GEN_1489); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1492 = 8'hd5 == _GEN_1064 ? $signed(-16'shc9) : $signed(_GEN_1490); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1493 = 8'hd6 == _GEN_1064 ? $signed(-16'sh3ffb) : $signed(_GEN_1491); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1494 = 8'hd6 == _GEN_1064 ? $signed(16'sh192) : $signed(_GEN_1492); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1495 = 8'hd7 == _GEN_1064 ? $signed(-16'sh3fe1) : $signed(_GEN_1493); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1496 = 8'hd7 == _GEN_1064 ? $signed(16'sh3ed) : $signed(_GEN_1494); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1497 = 8'hd8 == _GEN_1064 ? $signed(-16'sh3fb1) : $signed(_GEN_1495); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1498 = 8'hd8 == _GEN_1064 ? $signed(16'sh646) : $signed(_GEN_1496); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1499 = 8'hd9 == _GEN_1064 ? $signed(-16'sh3f6b) : $signed(_GEN_1497); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1500 = 8'hd9 == _GEN_1064 ? $signed(16'sh89d) : $signed(_GEN_1498); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1501 = 8'hda == _GEN_1064 ? $signed(-16'sh3f0f) : $signed(_GEN_1499); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1502 = 8'hda == _GEN_1064 ? $signed(16'shaf1) : $signed(_GEN_1500); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1503 = 8'hdb == _GEN_1064 ? $signed(-16'sh3e9d) : $signed(_GEN_1501); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1504 = 8'hdb == _GEN_1064 ? $signed(16'shd41) : $signed(_GEN_1502); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1505 = 8'hdc == _GEN_1064 ? $signed(-16'sh3e15) : $signed(_GEN_1503); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1506 = 8'hdc == _GEN_1064 ? $signed(16'shf8d) : $signed(_GEN_1504); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1507 = 8'hdd == _GEN_1064 ? $signed(-16'sh3d78) : $signed(_GEN_1505); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1508 = 8'hdd == _GEN_1064 ? $signed(16'sh11d3) : $signed(_GEN_1506); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1509 = 8'hde == _GEN_1064 ? $signed(-16'sh3cc5) : $signed(_GEN_1507); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1510 = 8'hde == _GEN_1064 ? $signed(16'sh1413) : $signed(_GEN_1508); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1511 = 8'hdf == _GEN_1064 ? $signed(-16'sh3bfd) : $signed(_GEN_1509); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1512 = 8'hdf == _GEN_1064 ? $signed(16'sh164c) : $signed(_GEN_1510); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1513 = 8'he0 == _GEN_1064 ? $signed(-16'sh3b21) : $signed(_GEN_1511); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1514 = 8'he0 == _GEN_1064 ? $signed(16'sh187e) : $signed(_GEN_1512); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1515 = 8'he1 == _GEN_1064 ? $signed(-16'sh3a30) : $signed(_GEN_1513); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1516 = 8'he1 == _GEN_1064 ? $signed(16'sh1aa7) : $signed(_GEN_1514); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1517 = 8'he2 == _GEN_1064 ? $signed(-16'sh392b) : $signed(_GEN_1515); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1518 = 8'he2 == _GEN_1064 ? $signed(16'sh1cc6) : $signed(_GEN_1516); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1519 = 8'he3 == _GEN_1064 ? $signed(-16'sh3812) : $signed(_GEN_1517); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1520 = 8'he3 == _GEN_1064 ? $signed(16'sh1edc) : $signed(_GEN_1518); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1521 = 8'he4 == _GEN_1064 ? $signed(-16'sh36e5) : $signed(_GEN_1519); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1522 = 8'he4 == _GEN_1064 ? $signed(16'sh20e7) : $signed(_GEN_1520); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1523 = 8'he5 == _GEN_1064 ? $signed(-16'sh35a5) : $signed(_GEN_1521); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1524 = 8'he5 == _GEN_1064 ? $signed(16'sh22e7) : $signed(_GEN_1522); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1525 = 8'he6 == _GEN_1064 ? $signed(-16'sh3453) : $signed(_GEN_1523); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1526 = 8'he6 == _GEN_1064 ? $signed(16'sh24da) : $signed(_GEN_1524); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1527 = 8'he7 == _GEN_1064 ? $signed(-16'sh32ef) : $signed(_GEN_1525); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1528 = 8'he7 == _GEN_1064 ? $signed(16'sh26c1) : $signed(_GEN_1526); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1529 = 8'he8 == _GEN_1064 ? $signed(-16'sh3179) : $signed(_GEN_1527); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1530 = 8'he8 == _GEN_1064 ? $signed(16'sh289a) : $signed(_GEN_1528); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1531 = 8'he9 == _GEN_1064 ? $signed(-16'sh2ff2) : $signed(_GEN_1529); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1532 = 8'he9 == _GEN_1064 ? $signed(16'sh2a65) : $signed(_GEN_1530); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1533 = 8'hea == _GEN_1064 ? $signed(-16'sh2e5a) : $signed(_GEN_1531); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1534 = 8'hea == _GEN_1064 ? $signed(16'sh2c21) : $signed(_GEN_1532); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1535 = 8'heb == _GEN_1064 ? $signed(-16'sh2cb2) : $signed(_GEN_1533); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1536 = 8'heb == _GEN_1064 ? $signed(16'sh2dcf) : $signed(_GEN_1534); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1537 = 8'hec == _GEN_1064 ? $signed(-16'sh2afb) : $signed(_GEN_1535); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1538 = 8'hec == _GEN_1064 ? $signed(16'sh2f6c) : $signed(_GEN_1536); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1539 = 8'hed == _GEN_1064 ? $signed(-16'sh2935) : $signed(_GEN_1537); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1540 = 8'hed == _GEN_1064 ? $signed(16'sh30f9) : $signed(_GEN_1538); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1541 = 8'hee == _GEN_1064 ? $signed(-16'sh2760) : $signed(_GEN_1539); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1542 = 8'hee == _GEN_1064 ? $signed(16'sh3274) : $signed(_GEN_1540); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1543 = 8'hef == _GEN_1064 ? $signed(-16'sh257e) : $signed(_GEN_1541); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1544 = 8'hef == _GEN_1064 ? $signed(16'sh33df) : $signed(_GEN_1542); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1545 = 8'hf0 == _GEN_1064 ? $signed(-16'sh238e) : $signed(_GEN_1543); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1546 = 8'hf0 == _GEN_1064 ? $signed(16'sh3537) : $signed(_GEN_1544); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1547 = 8'hf1 == _GEN_1064 ? $signed(-16'sh2193) : $signed(_GEN_1545); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1548 = 8'hf1 == _GEN_1064 ? $signed(16'sh367d) : $signed(_GEN_1546); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1549 = 8'hf2 == _GEN_1064 ? $signed(-16'sh1f8c) : $signed(_GEN_1547); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1550 = 8'hf2 == _GEN_1064 ? $signed(16'sh37b0) : $signed(_GEN_1548); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1551 = 8'hf3 == _GEN_1064 ? $signed(-16'sh1d79) : $signed(_GEN_1549); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1552 = 8'hf3 == _GEN_1064 ? $signed(16'sh38cf) : $signed(_GEN_1550); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1553 = 8'hf4 == _GEN_1064 ? $signed(-16'sh1b5d) : $signed(_GEN_1551); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1554 = 8'hf4 == _GEN_1064 ? $signed(16'sh39db) : $signed(_GEN_1552); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1555 = 8'hf5 == _GEN_1064 ? $signed(-16'sh1937) : $signed(_GEN_1553); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1556 = 8'hf5 == _GEN_1064 ? $signed(16'sh3ad3) : $signed(_GEN_1554); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1557 = 8'hf6 == _GEN_1064 ? $signed(-16'sh1709) : $signed(_GEN_1555); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1558 = 8'hf6 == _GEN_1064 ? $signed(16'sh3bb6) : $signed(_GEN_1556); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1559 = 8'hf7 == _GEN_1064 ? $signed(-16'sh14d2) : $signed(_GEN_1557); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1560 = 8'hf7 == _GEN_1064 ? $signed(16'sh3c85) : $signed(_GEN_1558); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1561 = 8'hf8 == _GEN_1064 ? $signed(-16'sh1294) : $signed(_GEN_1559); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1562 = 8'hf8 == _GEN_1064 ? $signed(16'sh3d3f) : $signed(_GEN_1560); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1563 = 8'hf9 == _GEN_1064 ? $signed(-16'sh1050) : $signed(_GEN_1561); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1564 = 8'hf9 == _GEN_1064 ? $signed(16'sh3de3) : $signed(_GEN_1562); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1565 = 8'hfa == _GEN_1064 ? $signed(-16'she06) : $signed(_GEN_1563); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1566 = 8'hfa == _GEN_1064 ? $signed(16'sh3e72) : $signed(_GEN_1564); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1567 = 8'hfb == _GEN_1064 ? $signed(-16'shbb7) : $signed(_GEN_1565); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1568 = 8'hfb == _GEN_1064 ? $signed(16'sh3eeb) : $signed(_GEN_1566); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1569 = 8'hfc == _GEN_1064 ? $signed(-16'sh964) : $signed(_GEN_1567); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1570 = 8'hfc == _GEN_1064 ? $signed(16'sh3f4f) : $signed(_GEN_1568); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1571 = 8'hfd == _GEN_1064 ? $signed(-16'sh70e) : $signed(_GEN_1569); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1572 = 8'hfd == _GEN_1064 ? $signed(16'sh3f9c) : $signed(_GEN_1570); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1573 = 8'hfe == _GEN_1064 ? $signed(-16'sh4b5) : $signed(_GEN_1571); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1574 = 8'hfe == _GEN_1064 ? $signed(16'sh3fd4) : $signed(_GEN_1572); // @[SDFChainRadix22.scala 291:27]
  assign _GEN_1575 = 8'hff == _GEN_1064 ? $signed(-16'sh25b) : $signed(_GEN_1573); // @[SDFChainRadix22.scala 291:27]
  assign twiddles_7_imag = 8'hff == _GEN_1064 ? $signed(16'sh3ff5) : $signed(_GEN_1574); // @[SDFChainRadix22.scala 291:27]
  assign _T_2096 = $signed(_GEN_1575) + $signed(twiddles_7_imag); // @[FixedPointTypeClass.scala 24:22]
  assign outputWires_6_real = sdf_stages_6_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign outputWires_6_imag = sdf_stages_6_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign _T_2097 = $signed(outputWires_6_real) + $signed(outputWires_6_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_2098 = $signed(outputWires_6_imag) - $signed(outputWires_6_real); // @[FixedPointTypeClass.scala 33:22]
  assign _GEN_2121 = {{1{outputWires_6_real[15]}},outputWires_6_real}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_2099 = $signed(_GEN_2121) * $signed(_T_2096); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2122 = {{1{twiddles_7_imag[15]}},twiddles_7_imag}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_2100 = $signed(_T_2097) * $signed(_GEN_2122); // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_2123 = {{1{_GEN_1575[15]}},_GEN_1575}; // @[FixedPointTypeClass.scala 211:35]
  assign _T_2101 = $signed(_T_2098) * $signed(_GEN_2123); // @[FixedPointTypeClass.scala 211:35]
  assign _T_2102 = $signed(_T_2099) - $signed(_T_2100); // @[FixedPointTypeClass.scala 33:22]
  assign _T_2103 = $signed(_T_2099) + $signed(_T_2101); // @[FixedPointTypeClass.scala 24:22]
  assign _T_2109 = $signed(_T_2102) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_2110 = _T_2109[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_2113 = $signed(_T_2103) + 34'sh2000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_2114 = _T_2113[33:14]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_2121 = sdf_stages_8_io_cntr < 9'h100; // @[SDFChainRadix22.scala 328:32]
  assign _T_2122 = sdf_stages_8_io_cntr < 9'h180; // @[SDFChainRadix22.scala 328:78]
  assign _T_2123 = _T_2122 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 328:65]
  assign _T_2124 = _T_2121 ? 1'h0 : _T_2123; // @[SDFChainRadix22.scala 328:19]
  assign outputWires_7_real = sdf_stages_7_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _T_2130 = 16'sh0 - $signed(outputWires_7_real); // @[FixedPointTypeClass.scala 39:43]
  assign outputWires_7_imag = sdf_stages_7_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 320:30]
  assign _GEN_2091 = 4'h1 == _T_48[3:0] ? $signed(outputWires_1_real) : $signed(outputWires_0_real); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2092 = 4'h1 == _T_48[3:0] ? $signed(outputWires_1_imag) : $signed(outputWires_0_imag); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2093 = 4'h2 == _T_48[3:0] ? $signed(outputWires_2_real) : $signed(_GEN_2091); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2094 = 4'h2 == _T_48[3:0] ? $signed(outputWires_2_imag) : $signed(_GEN_2092); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2095 = 4'h3 == _T_48[3:0] ? $signed(outputWires_3_real) : $signed(_GEN_2093); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2096 = 4'h3 == _T_48[3:0] ? $signed(outputWires_3_imag) : $signed(_GEN_2094); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2097 = 4'h4 == _T_48[3:0] ? $signed(outputWires_4_real) : $signed(_GEN_2095); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2098 = 4'h4 == _T_48[3:0] ? $signed(outputWires_4_imag) : $signed(_GEN_2096); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2099 = 4'h5 == _T_48[3:0] ? $signed(outputWires_5_real) : $signed(_GEN_2097); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2100 = 4'h5 == _T_48[3:0] ? $signed(outputWires_5_imag) : $signed(_GEN_2098); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2101 = 4'h6 == _T_48[3:0] ? $signed(outputWires_6_real) : $signed(_GEN_2099); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2102 = 4'h6 == _T_48[3:0] ? $signed(outputWires_6_imag) : $signed(_GEN_2100); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2103 = 4'h7 == _T_48[3:0] ? $signed(outputWires_7_real) : $signed(_GEN_2101); // @[SDFChainRadix22.scala 364:24]
  assign _GEN_2104 = 4'h7 == _T_48[3:0] ? $signed(outputWires_7_imag) : $signed(_GEN_2102); // @[SDFChainRadix22.scala 364:24]
  assign outputWires_8_real = sdf_stages_8_io_out_real; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign _GEN_2105 = 4'h8 == _T_48[3:0] ? $signed(outputWires_8_real) : $signed(_GEN_2103); // @[SDFChainRadix22.scala 364:24]
  assign outputWires_8_imag = sdf_stages_8_io_out_imag; // @[SDFChainRadix22.scala 43:111 SDFChainRadix22.scala 339:32]
  assign _GEN_2106 = 4'h8 == _T_48[3:0] ? $signed(outputWires_8_imag) : $signed(_GEN_2104); // @[SDFChainRadix22.scala 364:24]
  assign _T_2140 = ~initialOutDone; // @[SDFChainRadix22.scala 368:33]
  assign _T_2141 = state != 2'h2; // @[SDFChainRadix22.scala 368:127]
  assign _T_2142 = io_out_ready & _T_2141; // @[SDFChainRadix22.scala 368:117]
  assign _GEN_2124 = {$signed(_GEN_2106), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_2107 = {{2{_GEN_2124[29]}},_GEN_2124}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_2125 = {$signed(_GEN_2105), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_2108 = {{2{_GEN_2125[29]}},_GEN_2125}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_2126 = _GEN_2108[31:14]; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 396:27]
  assign _GEN_2128 = _GEN_2107[31:14]; // @[SDFChainRadix22.scala 63:26 SDFChainRadix22.scala 384:22 SDFChainRadix22.scala 397:27]
  assign io_in_ready = _T_2140 | _T_2142; // @[SDFChainRadix22.scala 368:15]
  assign io_out_valid = enableInit & initialOutDone; // @[SDFChainRadix22.scala 401:18]
  assign io_out_bits_real = _GEN_2126[15:0]; // @[SDFChainRadix22.scala 400:17]
  assign io_out_bits_imag = _GEN_2128[15:0]; // @[SDFChainRadix22.scala 400:17]
  assign io_lastOut = pktEnd & _T_83; // @[SDFChainRadix22.scala 428:14]
  assign io_busy = state != 2'h0; // @[SDFChainRadix22.scala 430:11]
  assign sdf_stages_0_clock = clock;
  assign sdf_stages_0_io_in_real = io_in_bits_real; // @[SDFChainRadix22.scala 347:23]
  assign sdf_stages_0_io_in_imag = io_in_bits_imag; // @[SDFChainRadix22.scala 347:23]
  assign sdf_stages_0_io_cntr = {{8'd0}, _T_166[0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_0_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_1_clock = clock;
  assign sdf_stages_1_io_in_real = _T_275[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_1_io_in_imag = _T_279[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_1_io_cntr = {{7'd0}, _T_173[1:0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_1_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_2_clock = clock;
  assign sdf_stages_2_io_in_real = _T_289 ? $signed(outputWires_1_imag) : $signed(outputWires_1_real); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_2_io_in_imag = _T_289 ? $signed(_T_295) : $signed(outputWires_1_imag); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_2_io_cntr = {{6'd0}, _T_180[2:0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_2_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_3_clock = clock;
  assign sdf_stages_3_io_in_real = _T_407[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_3_io_in_imag = _T_411[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_3_io_cntr = {{5'd0}, _T_187[3:0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_3_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_4_clock = clock;
  assign sdf_stages_4_io_in_real = _T_421 ? $signed(outputWires_3_imag) : $signed(outputWires_3_real); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_4_io_in_imag = _T_421 ? $signed(_T_427) : $signed(outputWires_3_imag); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_4_io_cntr = {{4'd0}, _T_194[4:0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_4_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_5_clock = clock;
  assign sdf_stages_5_io_in_real = _T_779[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_5_io_in_imag = _T_783[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_5_io_cntr = {{3'd0}, _T_201[5:0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_5_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_6_clock = clock;
  assign sdf_stages_6_io_in_real = _T_793 ? $signed(outputWires_5_imag) : $signed(outputWires_5_real); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_6_io_in_imag = _T_793 ? $signed(_T_799) : $signed(outputWires_5_imag); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_6_io_cntr = {{2'd0}, _T_208[6:0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_6_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_7_clock = clock;
  assign sdf_stages_7_io_in_real = _T_2110[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_7_io_in_imag = _T_2114[15:0]; // @[SDFChainRadix22.scala 319:21]
  assign sdf_stages_7_io_cntr = {{1'd0}, _T_215[7:0]}; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_7_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
  assign sdf_stages_8_clock = clock;
  assign sdf_stages_8_reset = reset;
  assign sdf_stages_8_io_in_real = _T_2124 ? $signed(outputWires_7_imag) : $signed(outputWires_7_real); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_8_io_in_imag = _T_2124 ? $signed(_T_2130) : $signed(outputWires_7_imag); // @[SDFChainRadix22.scala 340:23]
  assign sdf_stages_8_io_cntr = cntr_wires_0 - _T_220; // @[SDFChainRadix22.scala 224:16]
  assign sdf_stages_8_io_en = _T_46 | _T_122; // @[SDFChainRadix22.scala 223:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  initialOutDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cnt = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cntValidOut = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_53) begin
      if (_T_46) begin
        state <= 2'h1;
      end
    end else if (_T_56) begin
      if (fireLast) begin
        state <= 2'h2;
      end
    end else if (_T_57) begin
      if (io_lastOut) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      initialOutDone <= 1'h0;
    end else begin
      initialOutDone <= _GEN_46;
    end
    if (reset) begin
      cnt <= 10'h0;
    end else if (_T_62) begin
      cnt <= 10'h0;
    end else if (enableInit) begin
      cnt <= _T_125;
    end
    if (reset) begin
      cntValidOut <= 9'h0;
    end else if (_T_77) begin
      cntValidOut <= 9'h0;
    end else if (_T_61) begin
      cntValidOut <= _T_80;
    end
  end
endmodule
module SDFFFT_size_512_width_16_radix_22_bitreverse_0(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  output        io_lastOut,
  input         io_lastIn,
  output        io_busy
);
  wire  SDFChainRadix22_clock; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_reset; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_io_in_ready; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_io_in_valid; // @[SDFFFT.scala 219:119]
  wire [15:0] SDFChainRadix22_io_in_bits_real; // @[SDFFFT.scala 219:119]
  wire [15:0] SDFChainRadix22_io_in_bits_imag; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_io_out_ready; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_io_out_valid; // @[SDFFFT.scala 219:119]
  wire [15:0] SDFChainRadix22_io_out_bits_real; // @[SDFFFT.scala 219:119]
  wire [15:0] SDFChainRadix22_io_out_bits_imag; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_io_lastOut; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_io_lastIn; // @[SDFFFT.scala 219:119]
  wire  SDFChainRadix22_io_busy; // @[SDFFFT.scala 219:119]
  reg [8:0] cntWin; // @[SDFFFT.scala 71:23]
  reg [31:0] _RAND_0;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire [8:0] _T_6; // @[SDFFFT.scala 80:22]
  wire [8:0] _T_8; // @[SDFFFT.scala 82:44]
  wire  _T_9; // @[SDFFFT.scala 82:29]
  wire  _T_10; // @[SDFFFT.scala 82:19]
  wire [7:0] _T_85; // @[Bitwise.scala 103:31]
  wire [7:0] _T_87; // @[Bitwise.scala 103:65]
  wire [7:0] _T_89; // @[Bitwise.scala 103:75]
  wire [7:0] _T_90; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_522; // @[Bitwise.scala 103:31]
  wire [7:0] _T_95; // @[Bitwise.scala 103:31]
  wire [7:0] _T_97; // @[Bitwise.scala 103:65]
  wire [7:0] _T_99; // @[Bitwise.scala 103:75]
  wire [7:0] _T_100; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_523; // @[Bitwise.scala 103:31]
  wire [7:0] _T_105; // @[Bitwise.scala 103:31]
  wire [7:0] _T_107; // @[Bitwise.scala 103:65]
  wire [7:0] _T_109; // @[Bitwise.scala 103:75]
  wire [7:0] _T_110; // @[Bitwise.scala 103:39]
  wire [8:0] _T_143; // @[Cat.scala 29:58]
  wire [8:0] addrWin; // @[Mux.scala 87:16]
  wire [31:0] _T_152; // @[FixedPointTypeClass.scala 42:59]
  wire [31:0] _T_153; // @[FixedPointTypeClass.scala 42:59]
  wire [17:0] _GEN_526; // @[SDFFFT.scala 301:31 SDFFFT.scala 309:21]
  wire [17:0] _GEN_528; // @[SDFFFT.scala 302:31 SDFFFT.scala 309:21]
  SDFChainRadix22 SDFChainRadix22 ( // @[SDFFFT.scala 219:119]
    .clock(SDFChainRadix22_clock),
    .reset(SDFChainRadix22_reset),
    .io_in_ready(SDFChainRadix22_io_in_ready),
    .io_in_valid(SDFChainRadix22_io_in_valid),
    .io_in_bits_real(SDFChainRadix22_io_in_bits_real),
    .io_in_bits_imag(SDFChainRadix22_io_in_bits_imag),
    .io_out_ready(SDFChainRadix22_io_out_ready),
    .io_out_valid(SDFChainRadix22_io_out_valid),
    .io_out_bits_real(SDFChainRadix22_io_out_bits_real),
    .io_out_bits_imag(SDFChainRadix22_io_out_bits_imag),
    .io_lastOut(SDFChainRadix22_io_lastOut),
    .io_lastIn(SDFChainRadix22_io_lastIn),
    .io_busy(SDFChainRadix22_io_busy)
  );
  assign _T_4 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = cntWin + 9'h1; // @[SDFFFT.scala 80:22]
  assign _T_8 = 9'h0 - 9'h1; // @[SDFFFT.scala 82:44]
  assign _T_9 = cntWin == _T_8; // @[SDFFFT.scala 82:29]
  assign _T_10 = io_lastIn | _T_9; // @[SDFFFT.scala 82:19]
  assign _T_85 = {{4'd0}, cntWin[7:4]}; // @[Bitwise.scala 103:31]
  assign _T_87 = {cntWin[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_89 = _T_87 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_90 = _T_85 | _T_89; // @[Bitwise.scala 103:39]
  assign _GEN_522 = {{2'd0}, _T_90[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_95 = _GEN_522 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_97 = {_T_90[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_99 = _T_97 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_100 = _T_95 | _T_99; // @[Bitwise.scala 103:39]
  assign _GEN_523 = {{1'd0}, _T_100[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_105 = _GEN_523 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_107 = {_T_100[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_109 = _T_107 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_110 = _T_105 | _T_109; // @[Bitwise.scala 103:39]
  assign _T_143 = {_T_110,cntWin[8]}; // @[Cat.scala 29:58]
  assign addrWin = _T_143; // @[Mux.scala 87:16]
  assign _T_152 = $signed(io_in_bits_real) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  assign _T_153 = $signed(io_in_bits_imag) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  assign io_in_ready = SDFChainRadix22_io_in_ready; // @[SDFFFT.scala 305:23 SDFFFT.scala 309:21]
  assign io_out_valid = SDFChainRadix22_io_out_valid; // @[SDFFFT.scala 306:18 SDFFFT.scala 313:24]
  assign io_out_bits_real = SDFChainRadix22_io_out_bits_real; // @[SDFFFT.scala 306:18 SDFFFT.scala 311:23]
  assign io_out_bits_imag = SDFChainRadix22_io_out_bits_imag; // @[SDFFFT.scala 306:18 SDFFFT.scala 311:23]
  assign io_lastOut = SDFChainRadix22_io_lastOut; // @[SDFFFT.scala 317:20]
  assign io_busy = SDFChainRadix22_io_busy; // @[SDFFFT.scala 320:15]
  assign SDFChainRadix22_clock = clock;
  assign SDFChainRadix22_reset = reset;
  assign SDFChainRadix22_io_in_valid = io_in_valid; // @[SDFFFT.scala 304:27 SDFFFT.scala 309:21]
  assign _GEN_526 = _T_152[31:14]; // @[SDFFFT.scala 301:31 SDFFFT.scala 309:21]
  assign SDFChainRadix22_io_in_bits_real = _GEN_526[15:0]; // @[SDFFFT.scala 301:31 SDFFFT.scala 309:21]
  assign _GEN_528 = _T_153[31:14]; // @[SDFFFT.scala 302:31 SDFFFT.scala 309:21]
  assign SDFChainRadix22_io_in_bits_imag = _GEN_528[15:0]; // @[SDFFFT.scala 302:31 SDFFFT.scala 309:21]
  assign SDFChainRadix22_io_out_ready = io_out_ready; // @[SDFFFT.scala 306:18 SDFFFT.scala 314:28]
  assign SDFChainRadix22_io_lastIn = io_lastIn; // @[SDFFFT.scala 316:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cntWin = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cntWin <= 9'h0;
    end else if (_T_10) begin
      cntWin <= 9'h0;
    end else if (_T_4) begin
      cntWin <= _T_6;
    end
  end
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_extra,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_extra
);
  reg  _T_read [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_read__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_read__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_extra [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire  _T_extra__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_5;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_read__T_18_addr = value_1;
  assign _T_read__T_18_data = _T_read[_T_read__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_read__T_10_data = io_enq_bits_read;
  assign _T_read__T_10_addr = value;
  assign _T_read__T_10_mask = 1'h1;
  assign _T_read__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_extra__T_18_addr = value_1;
  assign _T_extra__T_18_data = _T_extra[_T_extra__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_extra__T_10_data = io_enq_bits_extra;
  assign _T_extra__T_10_addr = value;
  assign _T_extra__T_10_mask = 1'h1;
  assign _T_extra__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_read = _T_read__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_extra = _T_extra__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_read[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_extra[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_read__T_10_en & _T_read__T_10_mask) begin
      _T_read[_T_read__T_10_addr] <= _T_read__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_extra__T_10_en & _T_extra__T_10_mask) begin
      _T_extra[_T_extra__T_10_addr] <= _T_extra__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4FFTBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  fft_clock; // @[FFTBlock.scala 59:21]
  wire  fft_reset; // @[FFTBlock.scala 59:21]
  wire  fft_io_in_ready; // @[FFTBlock.scala 59:21]
  wire  fft_io_in_valid; // @[FFTBlock.scala 59:21]
  wire [15:0] fft_io_in_bits_real; // @[FFTBlock.scala 59:21]
  wire [15:0] fft_io_in_bits_imag; // @[FFTBlock.scala 59:21]
  wire  fft_io_out_ready; // @[FFTBlock.scala 59:21]
  wire  fft_io_out_valid; // @[FFTBlock.scala 59:21]
  wire [15:0] fft_io_out_bits_real; // @[FFTBlock.scala 59:21]
  wire [15:0] fft_io_out_bits_imag; // @[FFTBlock.scala 59:21]
  wire  fft_io_lastOut; // @[FFTBlock.scala 59:21]
  wire  fft_io_lastIn; // @[FFTBlock.scala 59:21]
  wire  fft_io_busy; // @[FFTBlock.scala 59:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  busy; // @[FFTBlock.scala 63:34]
  reg [31:0] _RAND_0;
  wire  _T_2; // @[RegisterRouter.scala 40:39]
  wire  _T_4; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_11; // @[RegisterRouter.scala 48:19]
  wire  _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_5; // @[RegisterRouter.scala 42:26]
  wire  _T_171; // @[RegisterRouter.scala 59:16]
  wire  _T_172_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_172_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_175; // @[RegisterRouter.scala 65:29]
  SDFFFT_size_512_width_16_radix_22_bitreverse_0 fft ( // @[FFTBlock.scala 59:21]
    .clock(fft_clock),
    .reset(fft_reset),
    .io_in_ready(fft_io_in_ready),
    .io_in_valid(fft_io_in_valid),
    .io_in_bits_real(fft_io_in_bits_real),
    .io_in_bits_imag(fft_io_in_bits_imag),
    .io_out_ready(fft_io_out_ready),
    .io_out_valid(fft_io_out_valid),
    .io_out_bits_real(fft_io_out_bits_real),
    .io_out_bits_imag(fft_io_out_bits_imag),
    .io_lastOut(fft_io_lastOut),
    .io_lastIn(fft_io_lastIn),
    .io_busy(fft_io_busy)
  );
  Queue_1 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_11[7:2] == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  assign _T_171 = _T_53 & busy; // @[RegisterRouter.scala 59:16]
  assign _T_172_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_172_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_175 = ~_T_172_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_172_valid & _T_175; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_172_valid & _T_172_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = fft_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = fft_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {fft_io_out_bits_real,fft_io_out_bits_imag}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = fft_io_lastOut; // @[LazyModule.scala 173:49]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_io_in_valid = auto_stream_in_valid; // @[FFTBlock.scala 124:24]
  assign fft_io_in_bits_real = auto_stream_in_bits_data[31:16]; // @[FFTBlock.scala 130:26]
  assign fft_io_in_bits_imag = auto_stream_in_bits_data[15:0]; // @[FFTBlock.scala 129:26]
  assign fft_io_out_ready = auto_stream_out_ready; // @[FFTBlock.scala 137:22]
  assign fft_io_lastIn = auto_stream_in_bits_last; // @[FFTBlock.scala 133:24]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_171}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_172_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      busy <= 1'h0;
    end else begin
      busy <= fft_io_busy;
    end
  end
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits
);
  reg [15:0] _T [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] _T__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12; // @[Counter.scala 39:22]
  wire [1:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_3(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
  reg  _T [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12; // @[Counter.scala 39:22]
  wire [1:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module MagJPLandSQRMagInst(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  input  [1:0]  io_sel,
  output        io_lastOut
);
  wire  Queue_clock; // @[Skid.scala 26:23]
  wire  Queue_reset; // @[Skid.scala 26:23]
  wire  Queue_io_enq_ready; // @[Skid.scala 26:23]
  wire  Queue_io_enq_valid; // @[Skid.scala 26:23]
  wire [15:0] Queue_io_enq_bits; // @[Skid.scala 26:23]
  wire  Queue_io_deq_ready; // @[Skid.scala 26:23]
  wire  Queue_io_deq_valid; // @[Skid.scala 26:23]
  wire [15:0] Queue_io_deq_bits; // @[Skid.scala 26:23]
  wire  Queue_1_clock; // @[Skid.scala 26:23]
  wire  Queue_1_reset; // @[Skid.scala 26:23]
  wire  Queue_1_io_enq_ready; // @[Skid.scala 26:23]
  wire  Queue_1_io_enq_valid; // @[Skid.scala 26:23]
  wire  Queue_1_io_enq_bits; // @[Skid.scala 26:23]
  wire  Queue_1_io_deq_ready; // @[Skid.scala 26:23]
  wire  Queue_1_io_deq_valid; // @[Skid.scala 26:23]
  wire  Queue_1_io_deq_bits; // @[Skid.scala 26:23]
  wire [15:0] _T_5; // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] absInReal; // @[FixedPointTypeClass.scala 247:8]
  wire [15:0] _T_9; // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] absInImag; // @[FixedPointTypeClass.scala 247:8]
  wire  _T_10; // @[FixedPointTypeClass.scala 55:59]
  wire [15:0] u; // @[Order.scala 56:31]
  wire  _T_11; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] v; // @[Order.scala 55:31]
  wire [12:0] _T_12; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] _GEN_16; // @[FixedPointTypeClass.scala 24:22]
  reg [16:0] _T_14; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [16:0] jplMagOp1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [12:0] _T_15; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] _GEN_17; // @[FixedPointTypeClass.scala 33:22]
  reg [16:0] tmpOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [14:0] _T_18; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  wire [16:0] _GEN_18; // @[FixedPointTypeClass.scala 24:22]
  reg [17:0] jplMagOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_21; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  wire [17:0] _T_22; // @[FixedPointTypeClass.scala 153:43]
  reg [31:0] _T_24; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  wire [17:0] _T_25; // @[FixedPointTypeClass.scala 153:43]
  reg [18:0] squared_magnitude; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  wire [21:0] _T_27; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [18:0] _T_29; // @[FixedPointTypeClass.scala 133:23]
  wire [18:0] _T_32; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] trim_squared_magnitude; // @[FixedPointTypeClass.scala 176:41]
  wire [17:0] _GEN_19; // @[FixedPointTypeClass.scala 55:59]
  wire  _T_33; // @[FixedPointTypeClass.scala 55:59]
  wire [17:0] jplMag; // @[Order.scala 56:31]
  reg [1:0] _T_34; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [1:0] _T_35; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  wire  _T_38; // @[Mux.scala 68:19]
  wire [18:0] _T_39; // @[Mux.scala 68:16]
  reg [1:0] queueCounter; // @[Skid.scala 27:31]
  reg [31:0] _RAND_10;
  wire  _T_48; // @[Skid.scala 35:31]
  wire  _T_49; // @[Skid.scala 35:68]
  wire  _T_50; // @[Skid.scala 35:89]
  wire  skidInData_ready; // @[Skid.scala 35:51]
  wire  _T_40; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_20; // @[Skid.scala 28:34]
  wire [2:0] _T_41; // @[Skid.scala 28:34]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_21; // @[Skid.scala 28:47]
  wire [3:0] _T_43; // @[Skid.scala 28:47]
  reg  _T_46; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg  _T_47; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  wire  _T_54; // @[Decoupled.scala 40:37]
  reg  _T_56; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg  _T_57; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [1:0] queueCounter_1; // @[Skid.scala 27:31]
  reg [31:0] _RAND_15;
  wire  _T_66; // @[Skid.scala 35:31]
  wire  _T_67; // @[Skid.scala 35:68]
  wire  _T_68; // @[Skid.scala 35:89]
  wire  _T_69; // @[Skid.scala 35:51]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_22; // @[Skid.scala 28:34]
  wire [2:0] _T_59; // @[Skid.scala 28:34]
  wire  _T_53_valid; // @[LogMagMuxTypes.scala 220:27 Skid.scala 37:15]
  wire  _T_60; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_23; // @[Skid.scala 28:47]
  wire [3:0] _T_61; // @[Skid.scala 28:47]
  reg  _T_64; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg  _T_65; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  Queue_2 Queue ( // @[Skid.scala 26:23]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_3 Queue_1 ( // @[Skid.scala 26:23]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  assign _T_5 = 16'sh0 - $signed(io_in_bits_real); // @[FixedPointTypeClass.scala 30:68]
  assign absInReal = io_in_bits_real[15] ? $signed(_T_5) : $signed(io_in_bits_real); // @[FixedPointTypeClass.scala 247:8]
  assign _T_9 = 16'sh0 - $signed(io_in_bits_imag); // @[FixedPointTypeClass.scala 30:68]
  assign absInImag = io_in_bits_imag[15] ? $signed(_T_9) : $signed(io_in_bits_imag); // @[FixedPointTypeClass.scala 247:8]
  assign _T_10 = $signed(absInReal) > $signed(absInImag); // @[FixedPointTypeClass.scala 55:59]
  assign u = _T_10 ? $signed(absInReal) : $signed(absInImag); // @[Order.scala 56:31]
  assign _T_11 = $signed(absInReal) < $signed(absInImag); // @[FixedPointTypeClass.scala 53:59]
  assign v = _T_11 ? $signed(absInReal) : $signed(absInImag); // @[Order.scala 55:31]
  assign _T_12 = v[15:3]; // @[FixedPointTypeClass.scala 117:50]
  assign _GEN_16 = {{3{_T_12[12]}},_T_12}; // @[FixedPointTypeClass.scala 24:22]
  assign _T_15 = u[15:3]; // @[FixedPointTypeClass.scala 117:50]
  assign _GEN_17 = {{3{_T_15[12]}},_T_15}; // @[FixedPointTypeClass.scala 33:22]
  assign _GEN_18 = {{2{_T_18[14]}},_T_18}; // @[FixedPointTypeClass.scala 24:22]
  assign _T_22 = _T_21[31:14]; // @[FixedPointTypeClass.scala 153:43]
  assign _T_25 = _T_24[31:14]; // @[FixedPointTypeClass.scala 153:43]
  assign _T_27 = {$signed(squared_magnitude), 3'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_29 = _T_27[21:3]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_32 = $signed(_T_29) + 19'sh4; // @[FixedPointTypeClass.scala 20:58]
  assign trim_squared_magnitude = _T_32[18:3]; // @[FixedPointTypeClass.scala 176:41]
  assign _GEN_19 = {{1{jplMagOp1[16]}},jplMagOp1}; // @[FixedPointTypeClass.scala 55:59]
  assign _T_33 = $signed(_GEN_19) > $signed(jplMagOp2); // @[FixedPointTypeClass.scala 55:59]
  assign jplMag = _T_33 ? $signed({{1{jplMagOp1[16]}},jplMagOp1}) : $signed(jplMagOp2); // @[Order.scala 56:31]
  assign _T_38 = 2'h0 == _T_35; // @[Mux.scala 68:19]
  assign _T_39 = _T_38 ? $signed(squared_magnitude) : $signed({{1{jplMag[17]}},jplMag}); // @[Mux.scala 68:16]
  assign _T_48 = queueCounter < 2'h3; // @[Skid.scala 35:31]
  assign _T_49 = queueCounter == 2'h3; // @[Skid.scala 35:68]
  assign _T_50 = _T_49 & io_out_ready; // @[Skid.scala 35:89]
  assign skidInData_ready = _T_48 | _T_50; // @[Skid.scala 35:51]
  assign _T_40 = skidInData_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = {{1'd0}, _T_40}; // @[Skid.scala 28:34]
  assign _T_41 = queueCounter + _GEN_20; // @[Skid.scala 28:34]
  assign _T_42 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = {{2'd0}, _T_42}; // @[Skid.scala 28:47]
  assign _T_43 = _T_41 - _GEN_21; // @[Skid.scala 28:47]
  assign _T_54 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_66 = queueCounter_1 < 2'h3; // @[Skid.scala 35:31]
  assign _T_67 = queueCounter_1 == 2'h3; // @[Skid.scala 35:68]
  assign _T_68 = _T_67 & io_out_ready; // @[Skid.scala 35:89]
  assign _T_69 = _T_66 | _T_68; // @[Skid.scala 35:51]
  assign _T_58 = _T_69 & io_in_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = {{1'd0}, _T_58}; // @[Skid.scala 28:34]
  assign _T_59 = queueCounter_1 + _GEN_22; // @[Skid.scala 28:34]
  assign _T_53_valid = Queue_1_io_deq_valid; // @[LogMagMuxTypes.scala 220:27 Skid.scala 37:15]
  assign _T_60 = io_out_ready & _T_53_valid; // @[Decoupled.scala 40:37]
  assign _GEN_23 = {{2'd0}, _T_60}; // @[Skid.scala 28:47]
  assign _T_61 = _T_59 - _GEN_23; // @[Skid.scala 28:47]
  assign io_in_ready = _T_48 | _T_50; // @[LogMagMuxTypes.scala 215:15]
  assign io_out_valid = Queue_io_deq_valid; // @[Skid.scala 37:15]
  assign io_out_bits = Queue_io_deq_bits; // @[Skid.scala 38:14]
  assign io_lastOut = Queue_1_io_deq_bits; // @[LogMagMuxTypes.scala 225:20]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_47; // @[Skid.scala 30:24]
  assign Queue_io_enq_bits = _T_39[15:0]; // @[LogMagMuxTypes.scala 216:37]
  assign Queue_io_deq_ready = io_out_ready; // @[Skid.scala 36:24]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_65; // @[Skid.scala 30:24]
  assign Queue_1_io_enq_bits = _T_57; // @[LogMagMuxTypes.scala 224:44]
  assign Queue_1_io_deq_ready = io_out_ready; // @[Skid.scala 36:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  jplMagOp1 = _RAND_1[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tmpOp2 = _RAND_2[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  jplMagOp2 = _RAND_4[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_24 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  squared_magnitude = _RAND_7[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_34 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_35 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  queueCounter = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_46 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_47 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_56 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_57 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  queueCounter_1 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_64 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_65 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= $signed(u) + $signed(_GEN_16);
    jplMagOp1 <= _T_14;
    tmpOp2 <= $signed(u) - $signed(_GEN_17);
    _T_18 <= v[15:1];
    jplMagOp2 <= $signed(tmpOp2) + $signed(_GEN_18);
    _T_21 <= $signed(absInReal) * $signed(absInReal);
    _T_24 <= $signed(absInImag) * $signed(absInImag);
    squared_magnitude <= $signed(_T_22) + $signed(_T_25);
    _T_34 <= io_sel;
    _T_35 <= _T_34;
    if (reset) begin
      queueCounter <= 2'h0;
    end else begin
      queueCounter <= _T_43[1:0];
    end
    if (reset) begin
      _T_46 <= 1'h0;
    end else begin
      _T_46 <= _T_40;
    end
    if (reset) begin
      _T_47 <= 1'h0;
    end else begin
      _T_47 <= _T_46;
    end
    _T_56 <= io_lastIn & _T_54;
    _T_57 <= _T_56;
    if (reset) begin
      queueCounter_1 <= 2'h0;
    end else begin
      queueCounter_1 <= _T_61[1:0];
    end
    if (reset) begin
      _T_64 <= 1'h0;
    end else begin
      _T_64 <= _T_58;
    end
    if (reset) begin
      _T_65 <= 1'h0;
    end else begin
      _T_65 <= _T_64;
    end
  end
endmodule
module LogMagMuxGenerator(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  input  [1:0]  io_sel,
  output        io_lastOut
);
  wire  magModule_clock; // @[LogMagMuxGenerator.scala 60:35]
  wire  magModule_reset; // @[LogMagMuxGenerator.scala 60:35]
  wire  magModule_io_in_ready; // @[LogMagMuxGenerator.scala 60:35]
  wire  magModule_io_in_valid; // @[LogMagMuxGenerator.scala 60:35]
  wire [15:0] magModule_io_in_bits_real; // @[LogMagMuxGenerator.scala 60:35]
  wire [15:0] magModule_io_in_bits_imag; // @[LogMagMuxGenerator.scala 60:35]
  wire  magModule_io_lastIn; // @[LogMagMuxGenerator.scala 60:35]
  wire  magModule_io_out_ready; // @[LogMagMuxGenerator.scala 60:35]
  wire  magModule_io_out_valid; // @[LogMagMuxGenerator.scala 60:35]
  wire [15:0] magModule_io_out_bits; // @[LogMagMuxGenerator.scala 60:35]
  wire [1:0] magModule_io_sel; // @[LogMagMuxGenerator.scala 60:35]
  wire  magModule_io_lastOut; // @[LogMagMuxGenerator.scala 60:35]
  MagJPLandSQRMagInst magModule ( // @[LogMagMuxGenerator.scala 60:35]
    .clock(magModule_clock),
    .reset(magModule_reset),
    .io_in_ready(magModule_io_in_ready),
    .io_in_valid(magModule_io_in_valid),
    .io_in_bits_real(magModule_io_in_bits_real),
    .io_in_bits_imag(magModule_io_in_bits_imag),
    .io_lastIn(magModule_io_lastIn),
    .io_out_ready(magModule_io_out_ready),
    .io_out_valid(magModule_io_out_valid),
    .io_out_bits(magModule_io_out_bits),
    .io_sel(magModule_io_sel),
    .io_lastOut(magModule_io_lastOut)
  );
  assign io_in_ready = magModule_io_in_ready; // @[LogMagMuxGenerator.scala 64:19]
  assign io_out_valid = magModule_io_out_valid; // @[LogMagMuxGenerator.scala 65:10]
  assign io_out_bits = magModule_io_out_bits; // @[LogMagMuxGenerator.scala 65:10]
  assign io_lastOut = magModule_io_lastOut; // @[LogMagMuxGenerator.scala 73:20]
  assign magModule_clock = clock;
  assign magModule_reset = reset;
  assign magModule_io_in_valid = io_in_valid; // @[LogMagMuxGenerator.scala 64:19]
  assign magModule_io_in_bits_real = io_in_bits_real; // @[LogMagMuxGenerator.scala 64:19]
  assign magModule_io_in_bits_imag = io_in_bits_imag; // @[LogMagMuxGenerator.scala 64:19]
  assign magModule_io_lastIn = io_lastIn; // @[LogMagMuxGenerator.scala 72:29]
  assign magModule_io_out_ready = io_out_ready; // @[LogMagMuxGenerator.scala 65:10]
  assign magModule_io_sel = io_sel; // @[LogMagMuxGenerator.scala 68:26]
endmodule
module AXI4LogMagMuxBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  input         auto_master_out_ready,
  output        auto_master_out_valid,
  output [15:0] auto_master_out_bits_data,
  output        auto_master_out_bits_last,
  output        auto_slave_in_ready,
  input         auto_slave_in_valid,
  input  [31:0] auto_slave_in_bits_data,
  input         auto_slave_in_bits_last
);
  wire  logMagMux_clock; // @[LogMagMuxDspBlock.scala 70:27]
  wire  logMagMux_reset; // @[LogMagMuxDspBlock.scala 70:27]
  wire  logMagMux_io_in_ready; // @[LogMagMuxDspBlock.scala 70:27]
  wire  logMagMux_io_in_valid; // @[LogMagMuxDspBlock.scala 70:27]
  wire [15:0] logMagMux_io_in_bits_real; // @[LogMagMuxDspBlock.scala 70:27]
  wire [15:0] logMagMux_io_in_bits_imag; // @[LogMagMuxDspBlock.scala 70:27]
  wire  logMagMux_io_lastIn; // @[LogMagMuxDspBlock.scala 70:27]
  wire  logMagMux_io_out_ready; // @[LogMagMuxDspBlock.scala 70:27]
  wire  logMagMux_io_out_valid; // @[LogMagMuxDspBlock.scala 70:27]
  wire [15:0] logMagMux_io_out_bits; // @[LogMagMuxDspBlock.scala 70:27]
  wire [1:0] logMagMux_io_sel; // @[LogMagMuxDspBlock.scala 70:27]
  wire  logMagMux_io_lastOut; // @[LogMagMuxDspBlock.scala 70:27]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  selReg; // @[LogMagMuxDspBlock.scala 75:25]
  reg [31:0] _RAND_0;
  wire  _T_2; // @[RegisterRouter.scala 40:39]
  wire  _T_3; // @[RegisterRouter.scala 40:26]
  wire  _T_4; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_11; // @[RegisterRouter.scala 48:19]
  wire  _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_5; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_14; // @[OneHot.scala 65:12]
  wire [1:0] _T_16; // @[Misc.scala 200:81]
  wire  _T_17; // @[Misc.scala 204:21]
  wire  _T_20; // @[Misc.scala 209:20]
  wire  _T_22; // @[Misc.scala 213:38]
  wire  _T_23; // @[Misc.scala 213:29]
  wire  _T_25; // @[Misc.scala 213:38]
  wire  _T_26; // @[Misc.scala 213:29]
  wire  _T_29; // @[Misc.scala 209:20]
  wire  _T_30; // @[Misc.scala 212:27]
  wire  _T_31; // @[Misc.scala 213:38]
  wire  _T_32; // @[Misc.scala 213:29]
  wire  _T_33; // @[Misc.scala 212:27]
  wire  _T_34; // @[Misc.scala 213:38]
  wire  _T_35; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 212:27]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_39; // @[Misc.scala 212:27]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire [3:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_63; // @[Bitwise.scala 72:12]
  wire [7:0] _T_65; // @[Bitwise.scala 72:12]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [31:0] _T_72; // @[Cat.scala 29:58]
  wire  _T_117; // @[RegisterRouter.scala 59:16]
  wire  _T_129; // @[RegisterRouter.scala 59:16]
  wire  _T_132; // @[RegisterRouter.scala 59:16]
  wire  _T_98; // @[RegisterRouter.scala 59:16]
  wire  _T_171; // @[RegisterRouter.scala 59:16]
  wire  _T_172_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_172_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_175; // @[RegisterRouter.scala 65:29]
  LogMagMuxGenerator logMagMux ( // @[LogMagMuxDspBlock.scala 70:27]
    .clock(logMagMux_clock),
    .reset(logMagMux_reset),
    .io_in_ready(logMagMux_io_in_ready),
    .io_in_valid(logMagMux_io_in_valid),
    .io_in_bits_real(logMagMux_io_in_bits_real),
    .io_in_bits_imag(logMagMux_io_in_bits_imag),
    .io_lastIn(logMagMux_io_lastIn),
    .io_out_ready(logMagMux_io_out_ready),
    .io_out_valid(logMagMux_io_out_valid),
    .io_out_bits(logMagMux_io_out_bits),
    .io_sel(logMagMux_io_sel),
    .io_lastOut(logMagMux_io_lastOut)
  );
  Queue_1 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_3 = auto_mem_in_ar_valid | _T_2; // @[RegisterRouter.scala 40:26]
  assign _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_11[7:2] == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  assign _T_14 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_16 = _T_14 | 2'h1; // @[Misc.scala 200:81]
  assign _T_17 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_20 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_22 = _T_16[1] & _T_20; // @[Misc.scala 213:38]
  assign _T_23 = _T_17 | _T_22; // @[Misc.scala 213:29]
  assign _T_25 = _T_16[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_26 = _T_17 | _T_25; // @[Misc.scala 213:29]
  assign _T_29 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_30 = _T_20 & _T_29; // @[Misc.scala 212:27]
  assign _T_31 = _T_16[0] & _T_30; // @[Misc.scala 213:38]
  assign _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  assign _T_33 = _T_20 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_34 = _T_16[0] & _T_33; // @[Misc.scala 213:38]
  assign _T_35 = _T_23 | _T_34; // @[Misc.scala 213:29]
  assign _T_36 = auto_mem_in_ar_bits_addr[1] & _T_29; // @[Misc.scala 212:27]
  assign _T_37 = _T_16[0] & _T_36; // @[Misc.scala 213:38]
  assign _T_38 = _T_26 | _T_37; // @[Misc.scala 213:29]
  assign _T_39 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_40 = _T_16[0] & _T_39; // @[Misc.scala 213:38]
  assign _T_41 = _T_26 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = {_T_41,_T_38,_T_35,_T_32}; // @[Cat.scala 29:58]
  assign _T_46 = auto_mem_in_ar_valid ? _T_44 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_63 = _T_46[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_65 = _T_46[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_67 = _T_46[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_46[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_72 = {_T_69,_T_67,_T_65,_T_63}; // @[Cat.scala 29:58]
  assign _T_117 = _T_3 & _T_47_ready; // @[RegisterRouter.scala 59:16]
  assign _T_129 = _T_117 & _T_4; // @[RegisterRouter.scala 59:16]
  assign _T_132 = _T_129 & _T_53; // @[RegisterRouter.scala 59:16]
  assign _T_98 = _T_132 & _T_72[0]; // @[RegisterRouter.scala 59:16]
  assign _T_171 = _T_53 & selReg; // @[RegisterRouter.scala 59:16]
  assign _T_172_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_172_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_175 = ~_T_172_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_172_valid & _T_175; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_172_valid & _T_172_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_master_out_valid = logMagMux_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_data = logMagMux_io_out_bits; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_last = logMagMux_io_lastOut; // @[LazyModule.scala 173:49]
  assign auto_slave_in_ready = logMagMux_io_in_ready; // @[LazyModule.scala 173:31]
  assign logMagMux_clock = clock;
  assign logMagMux_reset = reset;
  assign logMagMux_io_in_valid = auto_slave_in_valid; // @[LogMagMuxDspBlock.scala 87:30]
  assign logMagMux_io_in_bits_real = auto_slave_in_bits_data[31:16]; // @[LogMagMuxDspBlock.scala 88:30]
  assign logMagMux_io_in_bits_imag = auto_slave_in_bits_data[15:0]; // @[LogMagMuxDspBlock.scala 88:30]
  assign logMagMux_io_lastIn = auto_slave_in_bits_last; // @[LogMagMuxDspBlock.scala 91:31]
  assign logMagMux_io_out_ready = auto_master_out_ready; // @[LogMagMuxDspBlock.scala 96:28]
  assign logMagMux_io_sel = {{1'd0}, selReg}; // @[LogMagMuxDspBlock.scala 81:26]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_171}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_172_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  selReg = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      selReg <= 1'h0;
    end else if (_T_98) begin
      selReg <= auto_mem_in_w_bits_data[0];
    end
  end
endmodule
module AdjustableShiftRegisterStream(
  input         clock,
  input         reset,
  input  [6:0]  io_depth,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut,
  output [15:0] io_parallelOut_0,
  output [15:0] io_parallelOut_1,
  output [15:0] io_parallelOut_2,
  output [15:0] io_parallelOut_3,
  output [15:0] io_parallelOut_4,
  output [15:0] io_parallelOut_5,
  output [15:0] io_parallelOut_6,
  output [15:0] io_parallelOut_7,
  output [15:0] io_parallelOut_8,
  output [15:0] io_parallelOut_9,
  output [15:0] io_parallelOut_10,
  output [15:0] io_parallelOut_11,
  output [15:0] io_parallelOut_12,
  output [15:0] io_parallelOut_13,
  output [15:0] io_parallelOut_14,
  output [15:0] io_parallelOut_15,
  output [15:0] io_parallelOut_16,
  output [15:0] io_parallelOut_17,
  output [15:0] io_parallelOut_18,
  output [15:0] io_parallelOut_19,
  output [15:0] io_parallelOut_20,
  output [15:0] io_parallelOut_21,
  output [15:0] io_parallelOut_22,
  output [15:0] io_parallelOut_23,
  output [15:0] io_parallelOut_24,
  output [15:0] io_parallelOut_25,
  output [15:0] io_parallelOut_26,
  output [15:0] io_parallelOut_27,
  output [15:0] io_parallelOut_28,
  output [15:0] io_parallelOut_29,
  output [15:0] io_parallelOut_30,
  output [15:0] io_parallelOut_31,
  output [15:0] io_parallelOut_32,
  output [15:0] io_parallelOut_33,
  output [15:0] io_parallelOut_34,
  output [15:0] io_parallelOut_35,
  output [15:0] io_parallelOut_36,
  output [15:0] io_parallelOut_37,
  output [15:0] io_parallelOut_38,
  output [15:0] io_parallelOut_39,
  output [15:0] io_parallelOut_40,
  output [15:0] io_parallelOut_41,
  output [15:0] io_parallelOut_42,
  output [15:0] io_parallelOut_43,
  output [15:0] io_parallelOut_44,
  output [15:0] io_parallelOut_45,
  output [15:0] io_parallelOut_46,
  output [15:0] io_parallelOut_47,
  output [15:0] io_parallelOut_48,
  output [15:0] io_parallelOut_49,
  output [15:0] io_parallelOut_50,
  output [15:0] io_parallelOut_51,
  output [15:0] io_parallelOut_52,
  output [15:0] io_parallelOut_53,
  output [15:0] io_parallelOut_54,
  output [15:0] io_parallelOut_55,
  output [15:0] io_parallelOut_56,
  output [15:0] io_parallelOut_57,
  output [15:0] io_parallelOut_58,
  output [15:0] io_parallelOut_59,
  output [15:0] io_parallelOut_60,
  output [15:0] io_parallelOut_61,
  output [15:0] io_parallelOut_62,
  output [15:0] io_parallelOut_63,
  output [6:0]  io_cnt,
  output        io_regFull
);
  reg  InitialInDone; // @[CFARUtils.scala 379:30]
  reg [31:0] _RAND_0;
  reg  last; // @[CFARUtils.scala 380:21]
  reg [31:0] _RAND_1;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[CFARUtils.scala 385:34]
  wire  en; // @[CFARUtils.scala 385:25]
  wire  _T_3; // @[CFARUtils.scala 345:18]
  wire  _T_5; // @[CFARUtils.scala 345:11]
  wire  _T_6; // @[CFARUtils.scala 345:11]
  wire [6:0] _T_8; // @[CFARUtils.scala 350:87]
  wire  _T_9; // @[CFARUtils.scala 350:78]
  wire  _T_13; // @[CFARUtils.scala 350:78]
  wire  _T_14; // @[CFARUtils.scala 350:94]
  wire  _T_17; // @[CFARUtils.scala 350:78]
  wire  _T_18; // @[CFARUtils.scala 350:94]
  wire  _T_21; // @[CFARUtils.scala 350:78]
  wire  _T_22; // @[CFARUtils.scala 350:94]
  wire  _T_25; // @[CFARUtils.scala 350:78]
  wire  _T_26; // @[CFARUtils.scala 350:94]
  wire  _T_29; // @[CFARUtils.scala 350:78]
  wire  _T_30; // @[CFARUtils.scala 350:94]
  wire  _T_33; // @[CFARUtils.scala 350:78]
  wire  _T_34; // @[CFARUtils.scala 350:94]
  wire  _T_37; // @[CFARUtils.scala 350:78]
  wire  _T_38; // @[CFARUtils.scala 350:94]
  wire  _T_41; // @[CFARUtils.scala 350:78]
  wire  _T_42; // @[CFARUtils.scala 350:94]
  wire  _T_45; // @[CFARUtils.scala 350:78]
  wire  _T_46; // @[CFARUtils.scala 350:94]
  wire  _T_49; // @[CFARUtils.scala 350:78]
  wire  _T_50; // @[CFARUtils.scala 350:94]
  wire  _T_53; // @[CFARUtils.scala 350:78]
  wire  _T_54; // @[CFARUtils.scala 350:94]
  wire  _T_57; // @[CFARUtils.scala 350:78]
  wire  _T_58; // @[CFARUtils.scala 350:94]
  wire  _T_61; // @[CFARUtils.scala 350:78]
  wire  _T_62; // @[CFARUtils.scala 350:94]
  wire  _T_65; // @[CFARUtils.scala 350:78]
  wire  _T_66; // @[CFARUtils.scala 350:94]
  wire  _T_69; // @[CFARUtils.scala 350:78]
  wire  _T_70; // @[CFARUtils.scala 350:94]
  wire  _T_73; // @[CFARUtils.scala 350:78]
  wire  _T_74; // @[CFARUtils.scala 350:94]
  wire  _T_77; // @[CFARUtils.scala 350:78]
  wire  _T_78; // @[CFARUtils.scala 350:94]
  wire  _T_81; // @[CFARUtils.scala 350:78]
  wire  _T_82; // @[CFARUtils.scala 350:94]
  wire  _T_85; // @[CFARUtils.scala 350:78]
  wire  _T_86; // @[CFARUtils.scala 350:94]
  wire  _T_89; // @[CFARUtils.scala 350:78]
  wire  _T_90; // @[CFARUtils.scala 350:94]
  wire  _T_93; // @[CFARUtils.scala 350:78]
  wire  _T_94; // @[CFARUtils.scala 350:94]
  wire  _T_97; // @[CFARUtils.scala 350:78]
  wire  _T_98; // @[CFARUtils.scala 350:94]
  wire  _T_101; // @[CFARUtils.scala 350:78]
  wire  _T_102; // @[CFARUtils.scala 350:94]
  wire  _T_105; // @[CFARUtils.scala 350:78]
  wire  _T_106; // @[CFARUtils.scala 350:94]
  wire  _T_109; // @[CFARUtils.scala 350:78]
  wire  _T_110; // @[CFARUtils.scala 350:94]
  wire  _T_113; // @[CFARUtils.scala 350:78]
  wire  _T_114; // @[CFARUtils.scala 350:94]
  wire  _T_117; // @[CFARUtils.scala 350:78]
  wire  _T_118; // @[CFARUtils.scala 350:94]
  wire  _T_121; // @[CFARUtils.scala 350:78]
  wire  _T_122; // @[CFARUtils.scala 350:94]
  wire  _T_125; // @[CFARUtils.scala 350:78]
  wire  _T_126; // @[CFARUtils.scala 350:94]
  wire  _T_129; // @[CFARUtils.scala 350:78]
  wire  _T_130; // @[CFARUtils.scala 350:94]
  wire  _T_133; // @[CFARUtils.scala 350:78]
  wire  _T_134; // @[CFARUtils.scala 350:94]
  wire  _T_137; // @[CFARUtils.scala 350:78]
  wire  _T_138; // @[CFARUtils.scala 350:94]
  wire  _T_141; // @[CFARUtils.scala 350:78]
  wire  _T_142; // @[CFARUtils.scala 350:94]
  wire  _T_145; // @[CFARUtils.scala 350:78]
  wire  _T_146; // @[CFARUtils.scala 350:94]
  wire  _T_149; // @[CFARUtils.scala 350:78]
  wire  _T_150; // @[CFARUtils.scala 350:94]
  wire  _T_153; // @[CFARUtils.scala 350:78]
  wire  _T_154; // @[CFARUtils.scala 350:94]
  wire  _T_157; // @[CFARUtils.scala 350:78]
  wire  _T_158; // @[CFARUtils.scala 350:94]
  wire  _T_161; // @[CFARUtils.scala 350:78]
  wire  _T_162; // @[CFARUtils.scala 350:94]
  wire  _T_165; // @[CFARUtils.scala 350:78]
  wire  _T_166; // @[CFARUtils.scala 350:94]
  wire  _T_169; // @[CFARUtils.scala 350:78]
  wire  _T_170; // @[CFARUtils.scala 350:94]
  wire  _T_173; // @[CFARUtils.scala 350:78]
  wire  _T_174; // @[CFARUtils.scala 350:94]
  wire  _T_177; // @[CFARUtils.scala 350:78]
  wire  _T_178; // @[CFARUtils.scala 350:94]
  wire  _T_181; // @[CFARUtils.scala 350:78]
  wire  _T_182; // @[CFARUtils.scala 350:94]
  wire  _T_185; // @[CFARUtils.scala 350:78]
  wire  _T_186; // @[CFARUtils.scala 350:94]
  wire  _T_189; // @[CFARUtils.scala 350:78]
  wire  _T_190; // @[CFARUtils.scala 350:94]
  wire  _T_193; // @[CFARUtils.scala 350:78]
  wire  _T_194; // @[CFARUtils.scala 350:94]
  wire  _T_197; // @[CFARUtils.scala 350:78]
  wire  _T_198; // @[CFARUtils.scala 350:94]
  wire  _T_201; // @[CFARUtils.scala 350:78]
  wire  _T_202; // @[CFARUtils.scala 350:94]
  wire  _T_205; // @[CFARUtils.scala 350:78]
  wire  _T_206; // @[CFARUtils.scala 350:94]
  wire  _T_209; // @[CFARUtils.scala 350:78]
  wire  _T_210; // @[CFARUtils.scala 350:94]
  wire  _T_213; // @[CFARUtils.scala 350:78]
  wire  _T_214; // @[CFARUtils.scala 350:94]
  wire  _T_217; // @[CFARUtils.scala 350:78]
  wire  _T_218; // @[CFARUtils.scala 350:94]
  wire  _T_221; // @[CFARUtils.scala 350:78]
  wire  _T_222; // @[CFARUtils.scala 350:94]
  wire  _T_225; // @[CFARUtils.scala 350:78]
  wire  _T_226; // @[CFARUtils.scala 350:94]
  wire  _T_229; // @[CFARUtils.scala 350:78]
  wire  _T_230; // @[CFARUtils.scala 350:94]
  wire  _T_233; // @[CFARUtils.scala 350:78]
  wire  _T_234; // @[CFARUtils.scala 350:94]
  wire  _T_237; // @[CFARUtils.scala 350:78]
  wire  _T_238; // @[CFARUtils.scala 350:94]
  wire  _T_241; // @[CFARUtils.scala 350:78]
  wire  _T_242; // @[CFARUtils.scala 350:94]
  wire  _T_245; // @[CFARUtils.scala 350:78]
  wire  _T_246; // @[CFARUtils.scala 350:94]
  wire  _T_249; // @[CFARUtils.scala 350:78]
  wire  _T_250; // @[CFARUtils.scala 350:94]
  wire  _T_253; // @[CFARUtils.scala 350:78]
  wire  _T_254; // @[CFARUtils.scala 350:94]
  wire  _T_257; // @[CFARUtils.scala 350:78]
  wire  _T_258; // @[CFARUtils.scala 350:94]
  wire  _T_261; // @[CFARUtils.scala 350:78]
  wire  _T_262; // @[CFARUtils.scala 350:94]
  wire  activeRegs_63; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_263; // @[CFARUtils.scala 319:37]
  wire  activeRegs_62; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_264; // @[CFARUtils.scala 319:37]
  wire  activeRegs_61; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_265; // @[CFARUtils.scala 319:37]
  wire  activeRegs_60; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_266; // @[CFARUtils.scala 319:37]
  wire  activeRegs_59; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_267; // @[CFARUtils.scala 319:37]
  wire  activeRegs_58; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_268; // @[CFARUtils.scala 319:37]
  wire  activeRegs_57; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_269; // @[CFARUtils.scala 319:37]
  wire  activeRegs_56; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_270; // @[CFARUtils.scala 319:37]
  wire  activeRegs_55; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_271; // @[CFARUtils.scala 319:37]
  wire  activeRegs_54; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_272; // @[CFARUtils.scala 319:37]
  wire  activeRegs_53; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_273; // @[CFARUtils.scala 319:37]
  wire  activeRegs_52; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_274; // @[CFARUtils.scala 319:37]
  wire  activeRegs_51; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_275; // @[CFARUtils.scala 319:37]
  wire  activeRegs_50; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_276; // @[CFARUtils.scala 319:37]
  wire  activeRegs_49; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_277; // @[CFARUtils.scala 319:37]
  wire  activeRegs_48; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_278; // @[CFARUtils.scala 319:37]
  wire  activeRegs_47; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_279; // @[CFARUtils.scala 319:37]
  wire  activeRegs_46; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_280; // @[CFARUtils.scala 319:37]
  wire  activeRegs_45; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_281; // @[CFARUtils.scala 319:37]
  wire  activeRegs_44; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_282; // @[CFARUtils.scala 319:37]
  wire  activeRegs_43; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_283; // @[CFARUtils.scala 319:37]
  wire  activeRegs_42; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_284; // @[CFARUtils.scala 319:37]
  wire  activeRegs_41; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_285; // @[CFARUtils.scala 319:37]
  wire  activeRegs_40; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_286; // @[CFARUtils.scala 319:37]
  wire  activeRegs_39; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_287; // @[CFARUtils.scala 319:37]
  wire  activeRegs_38; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_288; // @[CFARUtils.scala 319:37]
  wire  activeRegs_37; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_289; // @[CFARUtils.scala 319:37]
  wire  activeRegs_36; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_290; // @[CFARUtils.scala 319:37]
  wire  activeRegs_35; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_291; // @[CFARUtils.scala 319:37]
  wire  activeRegs_34; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_292; // @[CFARUtils.scala 319:37]
  wire  activeRegs_33; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_293; // @[CFARUtils.scala 319:37]
  wire  activeRegs_32; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_294; // @[CFARUtils.scala 319:37]
  wire  activeRegs_31; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_295; // @[CFARUtils.scala 319:37]
  wire  activeRegs_30; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_296; // @[CFARUtils.scala 319:37]
  wire  activeRegs_29; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_297; // @[CFARUtils.scala 319:37]
  wire  activeRegs_28; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_298; // @[CFARUtils.scala 319:37]
  wire  activeRegs_27; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_299; // @[CFARUtils.scala 319:37]
  wire  activeRegs_26; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_300; // @[CFARUtils.scala 319:37]
  wire  activeRegs_25; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_301; // @[CFARUtils.scala 319:37]
  wire  activeRegs_24; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_302; // @[CFARUtils.scala 319:37]
  wire  activeRegs_23; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_303; // @[CFARUtils.scala 319:37]
  wire  activeRegs_22; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_304; // @[CFARUtils.scala 319:37]
  wire  activeRegs_21; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_305; // @[CFARUtils.scala 319:37]
  wire  activeRegs_20; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_306; // @[CFARUtils.scala 319:37]
  wire  activeRegs_19; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_307; // @[CFARUtils.scala 319:37]
  wire  activeRegs_18; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_308; // @[CFARUtils.scala 319:37]
  wire  activeRegs_17; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_309; // @[CFARUtils.scala 319:37]
  wire  activeRegs_16; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_310; // @[CFARUtils.scala 319:37]
  wire  activeRegs_15; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_311; // @[CFARUtils.scala 319:37]
  wire  activeRegs_14; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_312; // @[CFARUtils.scala 319:37]
  wire  activeRegs_13; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_313; // @[CFARUtils.scala 319:37]
  wire  activeRegs_12; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_314; // @[CFARUtils.scala 319:37]
  wire  activeRegs_11; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_315; // @[CFARUtils.scala 319:37]
  wire  activeRegs_10; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_316; // @[CFARUtils.scala 319:37]
  wire  activeRegs_9; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_317; // @[CFARUtils.scala 319:37]
  wire  activeRegs_8; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_318; // @[CFARUtils.scala 319:37]
  wire  activeRegs_7; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_319; // @[CFARUtils.scala 319:37]
  wire  activeRegs_6; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_320; // @[CFARUtils.scala 319:37]
  wire  activeRegs_5; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_321; // @[CFARUtils.scala 319:37]
  wire  activeRegs_4; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_322; // @[CFARUtils.scala 319:37]
  wire  activeRegs_3; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_323; // @[CFARUtils.scala 319:37]
  wire  activeRegs_2; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_324; // @[CFARUtils.scala 319:37]
  wire  activeRegs_1; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_325; // @[CFARUtils.scala 319:37]
  wire  activeRegs_0; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_326; // @[CFARUtils.scala 319:37]
  reg [15:0] adjShiftRegOut_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [15:0] adjShiftRegOut_1; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [15:0] adjShiftRegOut_2; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [15:0] adjShiftRegOut_3; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [15:0] adjShiftRegOut_4; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [15:0] adjShiftRegOut_5; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [15:0] adjShiftRegOut_6; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  reg [15:0] adjShiftRegOut_7; // @[Reg.scala 27:20]
  reg [31:0] _RAND_9;
  reg [15:0] adjShiftRegOut_8; // @[Reg.scala 27:20]
  reg [31:0] _RAND_10;
  reg [15:0] adjShiftRegOut_9; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg [15:0] adjShiftRegOut_10; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg [15:0] adjShiftRegOut_11; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg [15:0] adjShiftRegOut_12; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  reg [15:0] adjShiftRegOut_13; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  reg [15:0] adjShiftRegOut_14; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg [15:0] adjShiftRegOut_15; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  reg [15:0] adjShiftRegOut_16; // @[Reg.scala 27:20]
  reg [31:0] _RAND_18;
  reg [15:0] adjShiftRegOut_17; // @[Reg.scala 27:20]
  reg [31:0] _RAND_19;
  reg [15:0] adjShiftRegOut_18; // @[Reg.scala 27:20]
  reg [31:0] _RAND_20;
  reg [15:0] adjShiftRegOut_19; // @[Reg.scala 27:20]
  reg [31:0] _RAND_21;
  reg [15:0] adjShiftRegOut_20; // @[Reg.scala 27:20]
  reg [31:0] _RAND_22;
  reg [15:0] adjShiftRegOut_21; // @[Reg.scala 27:20]
  reg [31:0] _RAND_23;
  reg [15:0] adjShiftRegOut_22; // @[Reg.scala 27:20]
  reg [31:0] _RAND_24;
  reg [15:0] adjShiftRegOut_23; // @[Reg.scala 27:20]
  reg [31:0] _RAND_25;
  reg [15:0] adjShiftRegOut_24; // @[Reg.scala 27:20]
  reg [31:0] _RAND_26;
  reg [15:0] adjShiftRegOut_25; // @[Reg.scala 27:20]
  reg [31:0] _RAND_27;
  reg [15:0] adjShiftRegOut_26; // @[Reg.scala 27:20]
  reg [31:0] _RAND_28;
  reg [15:0] adjShiftRegOut_27; // @[Reg.scala 27:20]
  reg [31:0] _RAND_29;
  reg [15:0] adjShiftRegOut_28; // @[Reg.scala 27:20]
  reg [31:0] _RAND_30;
  reg [15:0] adjShiftRegOut_29; // @[Reg.scala 27:20]
  reg [31:0] _RAND_31;
  reg [15:0] adjShiftRegOut_30; // @[Reg.scala 27:20]
  reg [31:0] _RAND_32;
  reg [15:0] adjShiftRegOut_31; // @[Reg.scala 27:20]
  reg [31:0] _RAND_33;
  reg [15:0] adjShiftRegOut_32; // @[Reg.scala 27:20]
  reg [31:0] _RAND_34;
  reg [15:0] adjShiftRegOut_33; // @[Reg.scala 27:20]
  reg [31:0] _RAND_35;
  reg [15:0] adjShiftRegOut_34; // @[Reg.scala 27:20]
  reg [31:0] _RAND_36;
  reg [15:0] adjShiftRegOut_35; // @[Reg.scala 27:20]
  reg [31:0] _RAND_37;
  reg [15:0] adjShiftRegOut_36; // @[Reg.scala 27:20]
  reg [31:0] _RAND_38;
  reg [15:0] adjShiftRegOut_37; // @[Reg.scala 27:20]
  reg [31:0] _RAND_39;
  reg [15:0] adjShiftRegOut_38; // @[Reg.scala 27:20]
  reg [31:0] _RAND_40;
  reg [15:0] adjShiftRegOut_39; // @[Reg.scala 27:20]
  reg [31:0] _RAND_41;
  reg [15:0] adjShiftRegOut_40; // @[Reg.scala 27:20]
  reg [31:0] _RAND_42;
  reg [15:0] adjShiftRegOut_41; // @[Reg.scala 27:20]
  reg [31:0] _RAND_43;
  reg [15:0] adjShiftRegOut_42; // @[Reg.scala 27:20]
  reg [31:0] _RAND_44;
  reg [15:0] adjShiftRegOut_43; // @[Reg.scala 27:20]
  reg [31:0] _RAND_45;
  reg [15:0] adjShiftRegOut_44; // @[Reg.scala 27:20]
  reg [31:0] _RAND_46;
  reg [15:0] adjShiftRegOut_45; // @[Reg.scala 27:20]
  reg [31:0] _RAND_47;
  reg [15:0] adjShiftRegOut_46; // @[Reg.scala 27:20]
  reg [31:0] _RAND_48;
  reg [15:0] adjShiftRegOut_47; // @[Reg.scala 27:20]
  reg [31:0] _RAND_49;
  reg [15:0] adjShiftRegOut_48; // @[Reg.scala 27:20]
  reg [31:0] _RAND_50;
  reg [15:0] adjShiftRegOut_49; // @[Reg.scala 27:20]
  reg [31:0] _RAND_51;
  reg [15:0] adjShiftRegOut_50; // @[Reg.scala 27:20]
  reg [31:0] _RAND_52;
  reg [15:0] adjShiftRegOut_51; // @[Reg.scala 27:20]
  reg [31:0] _RAND_53;
  reg [15:0] adjShiftRegOut_52; // @[Reg.scala 27:20]
  reg [31:0] _RAND_54;
  reg [15:0] adjShiftRegOut_53; // @[Reg.scala 27:20]
  reg [31:0] _RAND_55;
  reg [15:0] adjShiftRegOut_54; // @[Reg.scala 27:20]
  reg [31:0] _RAND_56;
  reg [15:0] adjShiftRegOut_55; // @[Reg.scala 27:20]
  reg [31:0] _RAND_57;
  reg [15:0] adjShiftRegOut_56; // @[Reg.scala 27:20]
  reg [31:0] _RAND_58;
  reg [15:0] adjShiftRegOut_57; // @[Reg.scala 27:20]
  reg [31:0] _RAND_59;
  reg [15:0] adjShiftRegOut_58; // @[Reg.scala 27:20]
  reg [31:0] _RAND_60;
  reg [15:0] adjShiftRegOut_59; // @[Reg.scala 27:20]
  reg [31:0] _RAND_61;
  reg [15:0] adjShiftRegOut_60; // @[Reg.scala 27:20]
  reg [31:0] _RAND_62;
  reg [15:0] adjShiftRegOut_61; // @[Reg.scala 27:20]
  reg [31:0] _RAND_63;
  reg [15:0] adjShiftRegOut_62; // @[Reg.scala 27:20]
  reg [31:0] _RAND_64;
  reg [15:0] adjShiftRegOut_63; // @[Reg.scala 27:20]
  reg [31:0] _RAND_65;
  reg [6:0] cntIn; // @[CFARUtils.scala 390:23]
  reg [31:0] _RAND_66;
  wire  _T_395; // @[CFARUtils.scala 392:19]
  wire  _GEN_64; // @[CFARUtils.scala 392:36]
  wire [6:0] _T_398; // @[CFARUtils.scala 397:20]
  wire  _T_399; // @[CFARUtils.scala 400:18]
  wire  _T_402; // @[CFARUtils.scala 401:17]
  wire  _T_404; // @[CFARUtils.scala 401:36]
  wire  _GEN_66; // @[CFARUtils.scala 401:53]
  wire  _T_406; // @[CFARUtils.scala 406:36]
  wire  _T_407; // @[CFARUtils.scala 406:24]
  wire  _GEN_67; // @[CFARUtils.scala 406:45]
  wire  _T_409; // @[Decoupled.scala 40:37]
  wire  _T_672; // @[CFARUtils.scala 319:37]
  wire  _T_673; // @[CFARUtils.scala 319:37]
  wire  _T_674; // @[CFARUtils.scala 319:37]
  wire  _T_675; // @[CFARUtils.scala 319:37]
  wire  _T_676; // @[CFARUtils.scala 319:37]
  wire  _T_677; // @[CFARUtils.scala 319:37]
  wire  _T_678; // @[CFARUtils.scala 319:37]
  wire  _T_679; // @[CFARUtils.scala 319:37]
  wire  _T_680; // @[CFARUtils.scala 319:37]
  wire  _T_681; // @[CFARUtils.scala 319:37]
  wire  _T_682; // @[CFARUtils.scala 319:37]
  wire  _T_683; // @[CFARUtils.scala 319:37]
  wire  _T_684; // @[CFARUtils.scala 319:37]
  wire  _T_685; // @[CFARUtils.scala 319:37]
  wire  _T_686; // @[CFARUtils.scala 319:37]
  wire  _T_687; // @[CFARUtils.scala 319:37]
  wire  _T_688; // @[CFARUtils.scala 319:37]
  wire  _T_689; // @[CFARUtils.scala 319:37]
  wire  _T_690; // @[CFARUtils.scala 319:37]
  wire  _T_691; // @[CFARUtils.scala 319:37]
  wire  _T_692; // @[CFARUtils.scala 319:37]
  wire  _T_693; // @[CFARUtils.scala 319:37]
  wire  _T_694; // @[CFARUtils.scala 319:37]
  wire  _T_695; // @[CFARUtils.scala 319:37]
  wire  _T_696; // @[CFARUtils.scala 319:37]
  wire  _T_697; // @[CFARUtils.scala 319:37]
  wire  _T_698; // @[CFARUtils.scala 319:37]
  wire  _T_699; // @[CFARUtils.scala 319:37]
  wire  _T_700; // @[CFARUtils.scala 319:37]
  wire  _T_701; // @[CFARUtils.scala 319:37]
  wire  _T_702; // @[CFARUtils.scala 319:37]
  wire  _T_703; // @[CFARUtils.scala 319:37]
  wire  _T_704; // @[CFARUtils.scala 319:37]
  wire  _T_705; // @[CFARUtils.scala 319:37]
  wire  _T_706; // @[CFARUtils.scala 319:37]
  wire  _T_707; // @[CFARUtils.scala 319:37]
  wire  _T_708; // @[CFARUtils.scala 319:37]
  wire  _T_709; // @[CFARUtils.scala 319:37]
  wire  _T_710; // @[CFARUtils.scala 319:37]
  wire  _T_711; // @[CFARUtils.scala 319:37]
  wire  _T_712; // @[CFARUtils.scala 319:37]
  wire  _T_713; // @[CFARUtils.scala 319:37]
  wire  _T_714; // @[CFARUtils.scala 319:37]
  wire  _T_715; // @[CFARUtils.scala 319:37]
  wire  _T_716; // @[CFARUtils.scala 319:37]
  wire  _T_717; // @[CFARUtils.scala 319:37]
  wire  _T_718; // @[CFARUtils.scala 319:37]
  wire  _T_719; // @[CFARUtils.scala 319:37]
  wire  _T_720; // @[CFARUtils.scala 319:37]
  wire  _T_721; // @[CFARUtils.scala 319:37]
  wire  _T_722; // @[CFARUtils.scala 319:37]
  wire  _T_723; // @[CFARUtils.scala 319:37]
  wire  _T_724; // @[CFARUtils.scala 319:37]
  wire  _T_725; // @[CFARUtils.scala 319:37]
  wire  _T_726; // @[CFARUtils.scala 319:37]
  wire  _T_727; // @[CFARUtils.scala 319:37]
  wire  _T_728; // @[CFARUtils.scala 319:37]
  wire  _T_729; // @[CFARUtils.scala 319:37]
  wire  _T_730; // @[CFARUtils.scala 319:37]
  wire  _T_731; // @[CFARUtils.scala 319:37]
  wire  _T_732; // @[CFARUtils.scala 319:37]
  wire  _T_733; // @[CFARUtils.scala 319:37]
  wire  _T_734; // @[CFARUtils.scala 319:37]
  reg  _T_736; // @[Reg.scala 27:20]
  reg [31:0] _RAND_67;
  reg  _T_737; // @[Reg.scala 27:20]
  reg [31:0] _RAND_68;
  reg  _T_738; // @[Reg.scala 27:20]
  reg [31:0] _RAND_69;
  reg  _T_739; // @[Reg.scala 27:20]
  reg [31:0] _RAND_70;
  reg  _T_740; // @[Reg.scala 27:20]
  reg [31:0] _RAND_71;
  reg  _T_741; // @[Reg.scala 27:20]
  reg [31:0] _RAND_72;
  reg  _T_742; // @[Reg.scala 27:20]
  reg [31:0] _RAND_73;
  reg  _T_743; // @[Reg.scala 27:20]
  reg [31:0] _RAND_74;
  reg  _T_744; // @[Reg.scala 27:20]
  reg [31:0] _RAND_75;
  reg  _T_745; // @[Reg.scala 27:20]
  reg [31:0] _RAND_76;
  reg  _T_746; // @[Reg.scala 27:20]
  reg [31:0] _RAND_77;
  reg  _T_747; // @[Reg.scala 27:20]
  reg [31:0] _RAND_78;
  reg  _T_748; // @[Reg.scala 27:20]
  reg [31:0] _RAND_79;
  reg  _T_749; // @[Reg.scala 27:20]
  reg [31:0] _RAND_80;
  reg  _T_750; // @[Reg.scala 27:20]
  reg [31:0] _RAND_81;
  reg  _T_751; // @[Reg.scala 27:20]
  reg [31:0] _RAND_82;
  reg  _T_752; // @[Reg.scala 27:20]
  reg [31:0] _RAND_83;
  reg  _T_753; // @[Reg.scala 27:20]
  reg [31:0] _RAND_84;
  reg  _T_754; // @[Reg.scala 27:20]
  reg [31:0] _RAND_85;
  reg  _T_755; // @[Reg.scala 27:20]
  reg [31:0] _RAND_86;
  reg  _T_756; // @[Reg.scala 27:20]
  reg [31:0] _RAND_87;
  reg  _T_757; // @[Reg.scala 27:20]
  reg [31:0] _RAND_88;
  reg  _T_758; // @[Reg.scala 27:20]
  reg [31:0] _RAND_89;
  reg  _T_759; // @[Reg.scala 27:20]
  reg [31:0] _RAND_90;
  reg  _T_760; // @[Reg.scala 27:20]
  reg [31:0] _RAND_91;
  reg  _T_761; // @[Reg.scala 27:20]
  reg [31:0] _RAND_92;
  reg  _T_762; // @[Reg.scala 27:20]
  reg [31:0] _RAND_93;
  reg  _T_763; // @[Reg.scala 27:20]
  reg [31:0] _RAND_94;
  reg  _T_764; // @[Reg.scala 27:20]
  reg [31:0] _RAND_95;
  reg  _T_765; // @[Reg.scala 27:20]
  reg [31:0] _RAND_96;
  reg  _T_766; // @[Reg.scala 27:20]
  reg [31:0] _RAND_97;
  reg  _T_767; // @[Reg.scala 27:20]
  reg [31:0] _RAND_98;
  reg  _T_768; // @[Reg.scala 27:20]
  reg [31:0] _RAND_99;
  reg  _T_769; // @[Reg.scala 27:20]
  reg [31:0] _RAND_100;
  reg  _T_770; // @[Reg.scala 27:20]
  reg [31:0] _RAND_101;
  reg  _T_771; // @[Reg.scala 27:20]
  reg [31:0] _RAND_102;
  reg  _T_772; // @[Reg.scala 27:20]
  reg [31:0] _RAND_103;
  reg  _T_773; // @[Reg.scala 27:20]
  reg [31:0] _RAND_104;
  reg  _T_774; // @[Reg.scala 27:20]
  reg [31:0] _RAND_105;
  reg  _T_775; // @[Reg.scala 27:20]
  reg [31:0] _RAND_106;
  reg  _T_776; // @[Reg.scala 27:20]
  reg [31:0] _RAND_107;
  reg  _T_777; // @[Reg.scala 27:20]
  reg [31:0] _RAND_108;
  reg  _T_778; // @[Reg.scala 27:20]
  reg [31:0] _RAND_109;
  reg  _T_779; // @[Reg.scala 27:20]
  reg [31:0] _RAND_110;
  reg  _T_780; // @[Reg.scala 27:20]
  reg [31:0] _RAND_111;
  reg  _T_781; // @[Reg.scala 27:20]
  reg [31:0] _RAND_112;
  reg  _T_782; // @[Reg.scala 27:20]
  reg [31:0] _RAND_113;
  reg  _T_783; // @[Reg.scala 27:20]
  reg [31:0] _RAND_114;
  reg  _T_784; // @[Reg.scala 27:20]
  reg [31:0] _RAND_115;
  reg  _T_785; // @[Reg.scala 27:20]
  reg [31:0] _RAND_116;
  reg  _T_786; // @[Reg.scala 27:20]
  reg [31:0] _RAND_117;
  reg  _T_787; // @[Reg.scala 27:20]
  reg [31:0] _RAND_118;
  reg  _T_788; // @[Reg.scala 27:20]
  reg [31:0] _RAND_119;
  reg  _T_789; // @[Reg.scala 27:20]
  reg [31:0] _RAND_120;
  reg  _T_790; // @[Reg.scala 27:20]
  reg [31:0] _RAND_121;
  reg  _T_791; // @[Reg.scala 27:20]
  reg [31:0] _RAND_122;
  reg  _T_792; // @[Reg.scala 27:20]
  reg [31:0] _RAND_123;
  reg  _T_793; // @[Reg.scala 27:20]
  reg [31:0] _RAND_124;
  reg  _T_794; // @[Reg.scala 27:20]
  reg [31:0] _RAND_125;
  reg  _T_795; // @[Reg.scala 27:20]
  reg [31:0] _RAND_126;
  reg  _T_796; // @[Reg.scala 27:20]
  reg [31:0] _RAND_127;
  reg  _T_797; // @[Reg.scala 27:20]
  reg [31:0] _RAND_128;
  reg  _T_798; // @[Reg.scala 27:20]
  reg [31:0] _RAND_129;
  reg  _T_799; // @[Reg.scala 27:20]
  reg [31:0] _RAND_130;
  wire  _GEN_134; // @[CFARUtils.scala 414:17]
  wire  _GEN_135; // @[CFARUtils.scala 414:17]
  wire  _GEN_136; // @[CFARUtils.scala 414:17]
  wire  _GEN_137; // @[CFARUtils.scala 414:17]
  wire  _GEN_138; // @[CFARUtils.scala 414:17]
  wire  _GEN_139; // @[CFARUtils.scala 414:17]
  wire  _GEN_140; // @[CFARUtils.scala 414:17]
  wire  _GEN_141; // @[CFARUtils.scala 414:17]
  wire  _GEN_142; // @[CFARUtils.scala 414:17]
  wire  _GEN_143; // @[CFARUtils.scala 414:17]
  wire  _GEN_144; // @[CFARUtils.scala 414:17]
  wire  _GEN_145; // @[CFARUtils.scala 414:17]
  wire  _GEN_146; // @[CFARUtils.scala 414:17]
  wire  _GEN_147; // @[CFARUtils.scala 414:17]
  wire  _GEN_148; // @[CFARUtils.scala 414:17]
  wire  _GEN_149; // @[CFARUtils.scala 414:17]
  wire  _GEN_150; // @[CFARUtils.scala 414:17]
  wire  _GEN_151; // @[CFARUtils.scala 414:17]
  wire  _GEN_152; // @[CFARUtils.scala 414:17]
  wire  _GEN_153; // @[CFARUtils.scala 414:17]
  wire  _GEN_154; // @[CFARUtils.scala 414:17]
  wire  _GEN_155; // @[CFARUtils.scala 414:17]
  wire  _GEN_156; // @[CFARUtils.scala 414:17]
  wire  _GEN_157; // @[CFARUtils.scala 414:17]
  wire  _GEN_158; // @[CFARUtils.scala 414:17]
  wire  _GEN_159; // @[CFARUtils.scala 414:17]
  wire  _GEN_160; // @[CFARUtils.scala 414:17]
  wire  _GEN_161; // @[CFARUtils.scala 414:17]
  wire  _GEN_162; // @[CFARUtils.scala 414:17]
  wire  _GEN_163; // @[CFARUtils.scala 414:17]
  wire  _GEN_164; // @[CFARUtils.scala 414:17]
  wire  _GEN_165; // @[CFARUtils.scala 414:17]
  wire  _GEN_166; // @[CFARUtils.scala 414:17]
  wire  _GEN_167; // @[CFARUtils.scala 414:17]
  wire  _GEN_168; // @[CFARUtils.scala 414:17]
  wire  _GEN_169; // @[CFARUtils.scala 414:17]
  wire  _GEN_170; // @[CFARUtils.scala 414:17]
  wire  _GEN_171; // @[CFARUtils.scala 414:17]
  wire  _GEN_172; // @[CFARUtils.scala 414:17]
  wire  _GEN_173; // @[CFARUtils.scala 414:17]
  wire  _GEN_174; // @[CFARUtils.scala 414:17]
  wire  _GEN_175; // @[CFARUtils.scala 414:17]
  wire  _GEN_176; // @[CFARUtils.scala 414:17]
  wire  _GEN_177; // @[CFARUtils.scala 414:17]
  wire  _GEN_178; // @[CFARUtils.scala 414:17]
  wire  _GEN_179; // @[CFARUtils.scala 414:17]
  wire  _GEN_180; // @[CFARUtils.scala 414:17]
  wire  _GEN_181; // @[CFARUtils.scala 414:17]
  wire  _GEN_182; // @[CFARUtils.scala 414:17]
  wire  _GEN_183; // @[CFARUtils.scala 414:17]
  wire  _GEN_184; // @[CFARUtils.scala 414:17]
  wire  _GEN_185; // @[CFARUtils.scala 414:17]
  wire  _GEN_186; // @[CFARUtils.scala 414:17]
  wire  _GEN_187; // @[CFARUtils.scala 414:17]
  wire  _GEN_188; // @[CFARUtils.scala 414:17]
  wire  _GEN_189; // @[CFARUtils.scala 414:17]
  wire  _GEN_190; // @[CFARUtils.scala 414:17]
  wire  _GEN_191; // @[CFARUtils.scala 414:17]
  wire  _GEN_192; // @[CFARUtils.scala 414:17]
  wire  _GEN_193; // @[CFARUtils.scala 414:17]
  wire  _GEN_194; // @[CFARUtils.scala 414:17]
  wire  _GEN_195; // @[CFARUtils.scala 414:17]
  wire  _GEN_196; // @[CFARUtils.scala 414:17]
  wire  _T_804; // @[CFARUtils.scala 414:17]
  wire  _T_806; // @[CFARUtils.scala 420:36]
  wire  _T_808; // @[CFARUtils.scala 421:36]
  wire  _T_810; // @[CFARUtils.scala 426:37]
  wire  _T_813; // @[CFARUtils.scala 426:91]
  wire  _T_814; // @[CFARUtils.scala 426:75]
  wire [15:0] _GEN_201; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_202; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_203; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_204; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_205; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_206; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_207; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_208; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_209; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_210; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_211; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_212; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_213; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_214; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_215; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_216; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_217; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_218; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_219; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_220; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_221; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_222; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_223; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_224; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_225; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_226; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_227; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_228; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_229; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_230; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_231; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_232; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_233; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_234; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_235; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_236; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_237; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_238; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_239; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_240; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_241; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_242; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_243; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_244; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_245; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_246; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_247; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_248; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_249; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_250; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_251; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_252; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_253; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_254; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_255; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_256; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_257; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_258; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_259; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_260; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_261; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_262; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_263; // @[CFARUtils.scala 433:24]
  wire  _T_823; // @[CFARUtils.scala 436:70]
  wire  _T_824; // @[CFARUtils.scala 436:94]
  wire  _T_825; // @[CFARUtils.scala 436:85]
  assign _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = last & io_out_ready; // @[CFARUtils.scala 385:34]
  assign en = _T_1 | _T_2; // @[CFARUtils.scala 385:25]
  assign _T_3 = io_depth <= 7'h40; // @[CFARUtils.scala 345:18]
  assign _T_5 = _T_3 | reset; // @[CFARUtils.scala 345:11]
  assign _T_6 = ~_T_5; // @[CFARUtils.scala 345:11]
  assign _T_8 = io_depth - 7'h1; // @[CFARUtils.scala 350:87]
  assign _T_9 = 1'h1; // @[CFARUtils.scala 350:78]
  assign _T_13 = 7'h1 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_14 = _T_13; // @[CFARUtils.scala 350:94]
  assign _T_17 = 7'h2 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_18 = _T_17; // @[CFARUtils.scala 350:94]
  assign _T_21 = 7'h3 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_22 = _T_21; // @[CFARUtils.scala 350:94]
  assign _T_25 = 7'h4 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_26 = _T_25; // @[CFARUtils.scala 350:94]
  assign _T_29 = 7'h5 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_30 = _T_29; // @[CFARUtils.scala 350:94]
  assign _T_33 = 7'h6 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_34 = _T_33; // @[CFARUtils.scala 350:94]
  assign _T_37 = 7'h7 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_38 = _T_37; // @[CFARUtils.scala 350:94]
  assign _T_41 = 7'h8 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_42 = _T_41; // @[CFARUtils.scala 350:94]
  assign _T_45 = 7'h9 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_46 = _T_45; // @[CFARUtils.scala 350:94]
  assign _T_49 = 7'ha <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_50 = _T_49; // @[CFARUtils.scala 350:94]
  assign _T_53 = 7'hb <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_54 = _T_53; // @[CFARUtils.scala 350:94]
  assign _T_57 = 7'hc <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_58 = _T_57; // @[CFARUtils.scala 350:94]
  assign _T_61 = 7'hd <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_62 = _T_61; // @[CFARUtils.scala 350:94]
  assign _T_65 = 7'he <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_66 = _T_65; // @[CFARUtils.scala 350:94]
  assign _T_69 = 7'hf <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_70 = _T_69; // @[CFARUtils.scala 350:94]
  assign _T_73 = 7'h10 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_74 = _T_73; // @[CFARUtils.scala 350:94]
  assign _T_77 = 7'h11 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_78 = _T_77; // @[CFARUtils.scala 350:94]
  assign _T_81 = 7'h12 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_82 = _T_81; // @[CFARUtils.scala 350:94]
  assign _T_85 = 7'h13 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_86 = _T_85; // @[CFARUtils.scala 350:94]
  assign _T_89 = 7'h14 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_90 = _T_89; // @[CFARUtils.scala 350:94]
  assign _T_93 = 7'h15 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_94 = _T_93; // @[CFARUtils.scala 350:94]
  assign _T_97 = 7'h16 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_98 = _T_97; // @[CFARUtils.scala 350:94]
  assign _T_101 = 7'h17 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_102 = _T_101; // @[CFARUtils.scala 350:94]
  assign _T_105 = 7'h18 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_106 = _T_105; // @[CFARUtils.scala 350:94]
  assign _T_109 = 7'h19 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_110 = _T_109; // @[CFARUtils.scala 350:94]
  assign _T_113 = 7'h1a <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_114 = _T_113; // @[CFARUtils.scala 350:94]
  assign _T_117 = 7'h1b <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_118 = _T_117; // @[CFARUtils.scala 350:94]
  assign _T_121 = 7'h1c <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_122 = _T_121; // @[CFARUtils.scala 350:94]
  assign _T_125 = 7'h1d <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_126 = _T_125; // @[CFARUtils.scala 350:94]
  assign _T_129 = 7'h1e <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_130 = _T_129; // @[CFARUtils.scala 350:94]
  assign _T_133 = 7'h1f <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_134 = _T_133; // @[CFARUtils.scala 350:94]
  assign _T_137 = 7'h20 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_138 = _T_137; // @[CFARUtils.scala 350:94]
  assign _T_141 = 7'h21 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_142 = _T_141; // @[CFARUtils.scala 350:94]
  assign _T_145 = 7'h22 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_146 = _T_145; // @[CFARUtils.scala 350:94]
  assign _T_149 = 7'h23 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_150 = _T_149; // @[CFARUtils.scala 350:94]
  assign _T_153 = 7'h24 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_154 = _T_153; // @[CFARUtils.scala 350:94]
  assign _T_157 = 7'h25 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_158 = _T_157; // @[CFARUtils.scala 350:94]
  assign _T_161 = 7'h26 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_162 = _T_161; // @[CFARUtils.scala 350:94]
  assign _T_165 = 7'h27 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_166 = _T_165; // @[CFARUtils.scala 350:94]
  assign _T_169 = 7'h28 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_170 = _T_169; // @[CFARUtils.scala 350:94]
  assign _T_173 = 7'h29 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_174 = _T_173; // @[CFARUtils.scala 350:94]
  assign _T_177 = 7'h2a <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_178 = _T_177; // @[CFARUtils.scala 350:94]
  assign _T_181 = 7'h2b <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_182 = _T_181; // @[CFARUtils.scala 350:94]
  assign _T_185 = 7'h2c <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_186 = _T_185; // @[CFARUtils.scala 350:94]
  assign _T_189 = 7'h2d <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_190 = _T_189; // @[CFARUtils.scala 350:94]
  assign _T_193 = 7'h2e <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_194 = _T_193; // @[CFARUtils.scala 350:94]
  assign _T_197 = 7'h2f <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_198 = _T_197; // @[CFARUtils.scala 350:94]
  assign _T_201 = 7'h30 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_202 = _T_201; // @[CFARUtils.scala 350:94]
  assign _T_205 = 7'h31 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_206 = _T_205; // @[CFARUtils.scala 350:94]
  assign _T_209 = 7'h32 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_210 = _T_209; // @[CFARUtils.scala 350:94]
  assign _T_213 = 7'h33 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_214 = _T_213; // @[CFARUtils.scala 350:94]
  assign _T_217 = 7'h34 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_218 = _T_217; // @[CFARUtils.scala 350:94]
  assign _T_221 = 7'h35 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_222 = _T_221; // @[CFARUtils.scala 350:94]
  assign _T_225 = 7'h36 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_226 = _T_225; // @[CFARUtils.scala 350:94]
  assign _T_229 = 7'h37 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_230 = _T_229; // @[CFARUtils.scala 350:94]
  assign _T_233 = 7'h38 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_234 = _T_233; // @[CFARUtils.scala 350:94]
  assign _T_237 = 7'h39 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_238 = _T_237; // @[CFARUtils.scala 350:94]
  assign _T_241 = 7'h3a <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_242 = _T_241; // @[CFARUtils.scala 350:94]
  assign _T_245 = 7'h3b <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_246 = _T_245; // @[CFARUtils.scala 350:94]
  assign _T_249 = 7'h3c <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_250 = _T_249; // @[CFARUtils.scala 350:94]
  assign _T_253 = 7'h3d <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_254 = _T_253; // @[CFARUtils.scala 350:94]
  assign _T_257 = 7'h3e <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_258 = _T_257; // @[CFARUtils.scala 350:94]
  assign _T_261 = 7'h3f <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_262 = _T_261; // @[CFARUtils.scala 350:94]
  assign activeRegs_63 = _T_261; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_263 = _T_262 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_62 = _T_257; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_264 = _T_258 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_61 = _T_253; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_265 = _T_254 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_60 = _T_249; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_266 = _T_250 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_59 = _T_245; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_267 = _T_246 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_58 = _T_241; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_268 = _T_242 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_57 = _T_237; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_269 = _T_238 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_56 = _T_233; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_270 = _T_234 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_55 = _T_229; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_271 = _T_230 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_54 = _T_225; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_272 = _T_226 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_53 = _T_221; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_273 = _T_222 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_52 = _T_217; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_274 = _T_218 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_51 = _T_213; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_275 = _T_214 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_50 = _T_209; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_276 = _T_210 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_49 = _T_205; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_277 = _T_206 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_48 = _T_201; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_278 = _T_202 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_47 = _T_197; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_279 = _T_198 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_46 = _T_193; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_280 = _T_194 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_45 = _T_189; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_281 = _T_190 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_44 = _T_185; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_282 = _T_186 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_43 = _T_181; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_283 = _T_182 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_42 = _T_177; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_284 = _T_178 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_41 = _T_173; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_285 = _T_174 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_40 = _T_169; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_286 = _T_170 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_39 = _T_165; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_287 = _T_166 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_38 = _T_161; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_288 = _T_162 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_37 = _T_157; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_289 = _T_158 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_36 = _T_153; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_290 = _T_154 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_35 = _T_149; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_291 = _T_150 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_34 = _T_145; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_292 = _T_146 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_33 = _T_141; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_293 = _T_142 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_32 = _T_137; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_294 = _T_138 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_31 = _T_133; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_295 = _T_134 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_30 = _T_129; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_296 = _T_130 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_29 = _T_125; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_297 = _T_126 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_28 = _T_121; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_298 = _T_122 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_27 = _T_117; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_299 = _T_118 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_26 = _T_113; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_300 = _T_114 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_25 = _T_109; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_301 = _T_110 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_24 = _T_105; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_302 = _T_106 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_23 = _T_101; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_303 = _T_102 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_22 = _T_97; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_304 = _T_98 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_21 = _T_93; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_305 = _T_94 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_20 = _T_89; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_306 = _T_90 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_19 = _T_85; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_307 = _T_86 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_18 = _T_81; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_308 = _T_82 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_17 = _T_77; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_309 = _T_78 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_16 = _T_73; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_310 = _T_74 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_15 = _T_69; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_311 = _T_70 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_14 = _T_65; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_312 = _T_66 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_13 = _T_61; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_313 = _T_62 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_12 = _T_57; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_314 = _T_58 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_11 = _T_53; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_315 = _T_54 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_10 = _T_49; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_316 = _T_50 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_9 = _T_45; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_317 = _T_46 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_8 = _T_41; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_318 = _T_42 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_7 = _T_37; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_319 = _T_38 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_6 = _T_33; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_320 = _T_34 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_5 = _T_29; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_321 = _T_30 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_4 = _T_25; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_322 = _T_26 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_3 = _T_21; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_323 = _T_22 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_2 = _T_17; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_324 = _T_18 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_1 = _T_13; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_325 = _T_14 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_0 = 1'h1; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_326 = _T_9 & en; // @[CFARUtils.scala 319:37]
  assign _T_395 = io_lastIn & _T_1; // @[CFARUtils.scala 392:19]
  assign _GEN_64 = _T_395 | last; // @[CFARUtils.scala 392:36]
  assign _T_398 = cntIn + 7'h1; // @[CFARUtils.scala 397:20]
  assign _T_399 = io_depth > 7'h1; // @[CFARUtils.scala 400:18]
  assign _T_402 = cntIn == _T_8; // @[CFARUtils.scala 401:17]
  assign _T_404 = _T_402 & _T_1; // @[CFARUtils.scala 401:36]
  assign _GEN_66 = _T_404 | InitialInDone; // @[CFARUtils.scala 401:53]
  assign _T_406 = io_depth == 7'h1; // @[CFARUtils.scala 406:36]
  assign _T_407 = _T_1 & _T_406; // @[CFARUtils.scala 406:24]
  assign _GEN_67 = _T_407 | InitialInDone; // @[CFARUtils.scala 406:45]
  assign _T_409 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_672 = _T_261 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_673 = _T_257 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_674 = _T_253 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_675 = _T_249 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_676 = _T_245 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_677 = _T_241 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_678 = _T_237 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_679 = _T_233 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_680 = _T_229 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_681 = _T_225 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_682 = _T_221 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_683 = _T_217 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_684 = _T_213 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_685 = _T_209 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_686 = _T_205 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_687 = _T_201 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_688 = _T_197 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_689 = _T_193 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_690 = _T_189 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_691 = _T_185 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_692 = _T_181 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_693 = _T_177 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_694 = _T_173 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_695 = _T_169 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_696 = _T_165 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_697 = _T_161 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_698 = _T_157 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_699 = _T_153 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_700 = _T_149 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_701 = _T_145 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_702 = _T_141 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_703 = _T_137 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_704 = _T_133 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_705 = _T_129 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_706 = _T_125 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_707 = _T_121 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_708 = _T_117 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_709 = _T_113 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_710 = _T_109 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_711 = _T_105 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_712 = _T_101 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_713 = _T_97 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_714 = _T_93 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_715 = _T_89 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_716 = _T_85 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_717 = _T_81 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_718 = _T_77 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_719 = _T_73 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_720 = _T_69 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_721 = _T_65 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_722 = _T_61 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_723 = _T_57 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_724 = _T_53 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_725 = _T_49 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_726 = _T_45 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_727 = _T_41 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_728 = _T_37 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_729 = _T_33 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_730 = _T_29 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_731 = _T_25 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_732 = _T_21 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_733 = _T_17 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_734 = _T_13 & _T_409; // @[CFARUtils.scala 319:37]
  assign _GEN_134 = 6'h1 == _T_8[5:0] ? _T_737 : _T_736; // @[CFARUtils.scala 414:17]
  assign _GEN_135 = 6'h2 == _T_8[5:0] ? _T_738 : _GEN_134; // @[CFARUtils.scala 414:17]
  assign _GEN_136 = 6'h3 == _T_8[5:0] ? _T_739 : _GEN_135; // @[CFARUtils.scala 414:17]
  assign _GEN_137 = 6'h4 == _T_8[5:0] ? _T_740 : _GEN_136; // @[CFARUtils.scala 414:17]
  assign _GEN_138 = 6'h5 == _T_8[5:0] ? _T_741 : _GEN_137; // @[CFARUtils.scala 414:17]
  assign _GEN_139 = 6'h6 == _T_8[5:0] ? _T_742 : _GEN_138; // @[CFARUtils.scala 414:17]
  assign _GEN_140 = 6'h7 == _T_8[5:0] ? _T_743 : _GEN_139; // @[CFARUtils.scala 414:17]
  assign _GEN_141 = 6'h8 == _T_8[5:0] ? _T_744 : _GEN_140; // @[CFARUtils.scala 414:17]
  assign _GEN_142 = 6'h9 == _T_8[5:0] ? _T_745 : _GEN_141; // @[CFARUtils.scala 414:17]
  assign _GEN_143 = 6'ha == _T_8[5:0] ? _T_746 : _GEN_142; // @[CFARUtils.scala 414:17]
  assign _GEN_144 = 6'hb == _T_8[5:0] ? _T_747 : _GEN_143; // @[CFARUtils.scala 414:17]
  assign _GEN_145 = 6'hc == _T_8[5:0] ? _T_748 : _GEN_144; // @[CFARUtils.scala 414:17]
  assign _GEN_146 = 6'hd == _T_8[5:0] ? _T_749 : _GEN_145; // @[CFARUtils.scala 414:17]
  assign _GEN_147 = 6'he == _T_8[5:0] ? _T_750 : _GEN_146; // @[CFARUtils.scala 414:17]
  assign _GEN_148 = 6'hf == _T_8[5:0] ? _T_751 : _GEN_147; // @[CFARUtils.scala 414:17]
  assign _GEN_149 = 6'h10 == _T_8[5:0] ? _T_752 : _GEN_148; // @[CFARUtils.scala 414:17]
  assign _GEN_150 = 6'h11 == _T_8[5:0] ? _T_753 : _GEN_149; // @[CFARUtils.scala 414:17]
  assign _GEN_151 = 6'h12 == _T_8[5:0] ? _T_754 : _GEN_150; // @[CFARUtils.scala 414:17]
  assign _GEN_152 = 6'h13 == _T_8[5:0] ? _T_755 : _GEN_151; // @[CFARUtils.scala 414:17]
  assign _GEN_153 = 6'h14 == _T_8[5:0] ? _T_756 : _GEN_152; // @[CFARUtils.scala 414:17]
  assign _GEN_154 = 6'h15 == _T_8[5:0] ? _T_757 : _GEN_153; // @[CFARUtils.scala 414:17]
  assign _GEN_155 = 6'h16 == _T_8[5:0] ? _T_758 : _GEN_154; // @[CFARUtils.scala 414:17]
  assign _GEN_156 = 6'h17 == _T_8[5:0] ? _T_759 : _GEN_155; // @[CFARUtils.scala 414:17]
  assign _GEN_157 = 6'h18 == _T_8[5:0] ? _T_760 : _GEN_156; // @[CFARUtils.scala 414:17]
  assign _GEN_158 = 6'h19 == _T_8[5:0] ? _T_761 : _GEN_157; // @[CFARUtils.scala 414:17]
  assign _GEN_159 = 6'h1a == _T_8[5:0] ? _T_762 : _GEN_158; // @[CFARUtils.scala 414:17]
  assign _GEN_160 = 6'h1b == _T_8[5:0] ? _T_763 : _GEN_159; // @[CFARUtils.scala 414:17]
  assign _GEN_161 = 6'h1c == _T_8[5:0] ? _T_764 : _GEN_160; // @[CFARUtils.scala 414:17]
  assign _GEN_162 = 6'h1d == _T_8[5:0] ? _T_765 : _GEN_161; // @[CFARUtils.scala 414:17]
  assign _GEN_163 = 6'h1e == _T_8[5:0] ? _T_766 : _GEN_162; // @[CFARUtils.scala 414:17]
  assign _GEN_164 = 6'h1f == _T_8[5:0] ? _T_767 : _GEN_163; // @[CFARUtils.scala 414:17]
  assign _GEN_165 = 6'h20 == _T_8[5:0] ? _T_768 : _GEN_164; // @[CFARUtils.scala 414:17]
  assign _GEN_166 = 6'h21 == _T_8[5:0] ? _T_769 : _GEN_165; // @[CFARUtils.scala 414:17]
  assign _GEN_167 = 6'h22 == _T_8[5:0] ? _T_770 : _GEN_166; // @[CFARUtils.scala 414:17]
  assign _GEN_168 = 6'h23 == _T_8[5:0] ? _T_771 : _GEN_167; // @[CFARUtils.scala 414:17]
  assign _GEN_169 = 6'h24 == _T_8[5:0] ? _T_772 : _GEN_168; // @[CFARUtils.scala 414:17]
  assign _GEN_170 = 6'h25 == _T_8[5:0] ? _T_773 : _GEN_169; // @[CFARUtils.scala 414:17]
  assign _GEN_171 = 6'h26 == _T_8[5:0] ? _T_774 : _GEN_170; // @[CFARUtils.scala 414:17]
  assign _GEN_172 = 6'h27 == _T_8[5:0] ? _T_775 : _GEN_171; // @[CFARUtils.scala 414:17]
  assign _GEN_173 = 6'h28 == _T_8[5:0] ? _T_776 : _GEN_172; // @[CFARUtils.scala 414:17]
  assign _GEN_174 = 6'h29 == _T_8[5:0] ? _T_777 : _GEN_173; // @[CFARUtils.scala 414:17]
  assign _GEN_175 = 6'h2a == _T_8[5:0] ? _T_778 : _GEN_174; // @[CFARUtils.scala 414:17]
  assign _GEN_176 = 6'h2b == _T_8[5:0] ? _T_779 : _GEN_175; // @[CFARUtils.scala 414:17]
  assign _GEN_177 = 6'h2c == _T_8[5:0] ? _T_780 : _GEN_176; // @[CFARUtils.scala 414:17]
  assign _GEN_178 = 6'h2d == _T_8[5:0] ? _T_781 : _GEN_177; // @[CFARUtils.scala 414:17]
  assign _GEN_179 = 6'h2e == _T_8[5:0] ? _T_782 : _GEN_178; // @[CFARUtils.scala 414:17]
  assign _GEN_180 = 6'h2f == _T_8[5:0] ? _T_783 : _GEN_179; // @[CFARUtils.scala 414:17]
  assign _GEN_181 = 6'h30 == _T_8[5:0] ? _T_784 : _GEN_180; // @[CFARUtils.scala 414:17]
  assign _GEN_182 = 6'h31 == _T_8[5:0] ? _T_785 : _GEN_181; // @[CFARUtils.scala 414:17]
  assign _GEN_183 = 6'h32 == _T_8[5:0] ? _T_786 : _GEN_182; // @[CFARUtils.scala 414:17]
  assign _GEN_184 = 6'h33 == _T_8[5:0] ? _T_787 : _GEN_183; // @[CFARUtils.scala 414:17]
  assign _GEN_185 = 6'h34 == _T_8[5:0] ? _T_788 : _GEN_184; // @[CFARUtils.scala 414:17]
  assign _GEN_186 = 6'h35 == _T_8[5:0] ? _T_789 : _GEN_185; // @[CFARUtils.scala 414:17]
  assign _GEN_187 = 6'h36 == _T_8[5:0] ? _T_790 : _GEN_186; // @[CFARUtils.scala 414:17]
  assign _GEN_188 = 6'h37 == _T_8[5:0] ? _T_791 : _GEN_187; // @[CFARUtils.scala 414:17]
  assign _GEN_189 = 6'h38 == _T_8[5:0] ? _T_792 : _GEN_188; // @[CFARUtils.scala 414:17]
  assign _GEN_190 = 6'h39 == _T_8[5:0] ? _T_793 : _GEN_189; // @[CFARUtils.scala 414:17]
  assign _GEN_191 = 6'h3a == _T_8[5:0] ? _T_794 : _GEN_190; // @[CFARUtils.scala 414:17]
  assign _GEN_192 = 6'h3b == _T_8[5:0] ? _T_795 : _GEN_191; // @[CFARUtils.scala 414:17]
  assign _GEN_193 = 6'h3c == _T_8[5:0] ? _T_796 : _GEN_192; // @[CFARUtils.scala 414:17]
  assign _GEN_194 = 6'h3d == _T_8[5:0] ? _T_797 : _GEN_193; // @[CFARUtils.scala 414:17]
  assign _GEN_195 = 6'h3e == _T_8[5:0] ? _T_798 : _GEN_194; // @[CFARUtils.scala 414:17]
  assign _GEN_196 = 6'h3f == _T_8[5:0] ? _T_799 : _GEN_195; // @[CFARUtils.scala 414:17]
  assign _T_804 = _GEN_196 & _T_409; // @[CFARUtils.scala 414:17]
  assign _T_806 = ~InitialInDone; // @[CFARUtils.scala 420:36]
  assign _T_808 = ~last; // @[CFARUtils.scala 421:36]
  assign _T_810 = io_depth == 7'h0; // @[CFARUtils.scala 426:37]
  assign _T_813 = io_out_ready & _T_808; // @[CFARUtils.scala 426:91]
  assign _T_814 = _T_806 | _T_813; // @[CFARUtils.scala 426:75]
  assign _GEN_201 = 6'h1 == _T_8[5:0] ? $signed(adjShiftRegOut_1) : $signed(adjShiftRegOut_0); // @[CFARUtils.scala 433:24]
  assign _GEN_202 = 6'h2 == _T_8[5:0] ? $signed(adjShiftRegOut_2) : $signed(_GEN_201); // @[CFARUtils.scala 433:24]
  assign _GEN_203 = 6'h3 == _T_8[5:0] ? $signed(adjShiftRegOut_3) : $signed(_GEN_202); // @[CFARUtils.scala 433:24]
  assign _GEN_204 = 6'h4 == _T_8[5:0] ? $signed(adjShiftRegOut_4) : $signed(_GEN_203); // @[CFARUtils.scala 433:24]
  assign _GEN_205 = 6'h5 == _T_8[5:0] ? $signed(adjShiftRegOut_5) : $signed(_GEN_204); // @[CFARUtils.scala 433:24]
  assign _GEN_206 = 6'h6 == _T_8[5:0] ? $signed(adjShiftRegOut_6) : $signed(_GEN_205); // @[CFARUtils.scala 433:24]
  assign _GEN_207 = 6'h7 == _T_8[5:0] ? $signed(adjShiftRegOut_7) : $signed(_GEN_206); // @[CFARUtils.scala 433:24]
  assign _GEN_208 = 6'h8 == _T_8[5:0] ? $signed(adjShiftRegOut_8) : $signed(_GEN_207); // @[CFARUtils.scala 433:24]
  assign _GEN_209 = 6'h9 == _T_8[5:0] ? $signed(adjShiftRegOut_9) : $signed(_GEN_208); // @[CFARUtils.scala 433:24]
  assign _GEN_210 = 6'ha == _T_8[5:0] ? $signed(adjShiftRegOut_10) : $signed(_GEN_209); // @[CFARUtils.scala 433:24]
  assign _GEN_211 = 6'hb == _T_8[5:0] ? $signed(adjShiftRegOut_11) : $signed(_GEN_210); // @[CFARUtils.scala 433:24]
  assign _GEN_212 = 6'hc == _T_8[5:0] ? $signed(adjShiftRegOut_12) : $signed(_GEN_211); // @[CFARUtils.scala 433:24]
  assign _GEN_213 = 6'hd == _T_8[5:0] ? $signed(adjShiftRegOut_13) : $signed(_GEN_212); // @[CFARUtils.scala 433:24]
  assign _GEN_214 = 6'he == _T_8[5:0] ? $signed(adjShiftRegOut_14) : $signed(_GEN_213); // @[CFARUtils.scala 433:24]
  assign _GEN_215 = 6'hf == _T_8[5:0] ? $signed(adjShiftRegOut_15) : $signed(_GEN_214); // @[CFARUtils.scala 433:24]
  assign _GEN_216 = 6'h10 == _T_8[5:0] ? $signed(adjShiftRegOut_16) : $signed(_GEN_215); // @[CFARUtils.scala 433:24]
  assign _GEN_217 = 6'h11 == _T_8[5:0] ? $signed(adjShiftRegOut_17) : $signed(_GEN_216); // @[CFARUtils.scala 433:24]
  assign _GEN_218 = 6'h12 == _T_8[5:0] ? $signed(adjShiftRegOut_18) : $signed(_GEN_217); // @[CFARUtils.scala 433:24]
  assign _GEN_219 = 6'h13 == _T_8[5:0] ? $signed(adjShiftRegOut_19) : $signed(_GEN_218); // @[CFARUtils.scala 433:24]
  assign _GEN_220 = 6'h14 == _T_8[5:0] ? $signed(adjShiftRegOut_20) : $signed(_GEN_219); // @[CFARUtils.scala 433:24]
  assign _GEN_221 = 6'h15 == _T_8[5:0] ? $signed(adjShiftRegOut_21) : $signed(_GEN_220); // @[CFARUtils.scala 433:24]
  assign _GEN_222 = 6'h16 == _T_8[5:0] ? $signed(adjShiftRegOut_22) : $signed(_GEN_221); // @[CFARUtils.scala 433:24]
  assign _GEN_223 = 6'h17 == _T_8[5:0] ? $signed(adjShiftRegOut_23) : $signed(_GEN_222); // @[CFARUtils.scala 433:24]
  assign _GEN_224 = 6'h18 == _T_8[5:0] ? $signed(adjShiftRegOut_24) : $signed(_GEN_223); // @[CFARUtils.scala 433:24]
  assign _GEN_225 = 6'h19 == _T_8[5:0] ? $signed(adjShiftRegOut_25) : $signed(_GEN_224); // @[CFARUtils.scala 433:24]
  assign _GEN_226 = 6'h1a == _T_8[5:0] ? $signed(adjShiftRegOut_26) : $signed(_GEN_225); // @[CFARUtils.scala 433:24]
  assign _GEN_227 = 6'h1b == _T_8[5:0] ? $signed(adjShiftRegOut_27) : $signed(_GEN_226); // @[CFARUtils.scala 433:24]
  assign _GEN_228 = 6'h1c == _T_8[5:0] ? $signed(adjShiftRegOut_28) : $signed(_GEN_227); // @[CFARUtils.scala 433:24]
  assign _GEN_229 = 6'h1d == _T_8[5:0] ? $signed(adjShiftRegOut_29) : $signed(_GEN_228); // @[CFARUtils.scala 433:24]
  assign _GEN_230 = 6'h1e == _T_8[5:0] ? $signed(adjShiftRegOut_30) : $signed(_GEN_229); // @[CFARUtils.scala 433:24]
  assign _GEN_231 = 6'h1f == _T_8[5:0] ? $signed(adjShiftRegOut_31) : $signed(_GEN_230); // @[CFARUtils.scala 433:24]
  assign _GEN_232 = 6'h20 == _T_8[5:0] ? $signed(adjShiftRegOut_32) : $signed(_GEN_231); // @[CFARUtils.scala 433:24]
  assign _GEN_233 = 6'h21 == _T_8[5:0] ? $signed(adjShiftRegOut_33) : $signed(_GEN_232); // @[CFARUtils.scala 433:24]
  assign _GEN_234 = 6'h22 == _T_8[5:0] ? $signed(adjShiftRegOut_34) : $signed(_GEN_233); // @[CFARUtils.scala 433:24]
  assign _GEN_235 = 6'h23 == _T_8[5:0] ? $signed(adjShiftRegOut_35) : $signed(_GEN_234); // @[CFARUtils.scala 433:24]
  assign _GEN_236 = 6'h24 == _T_8[5:0] ? $signed(adjShiftRegOut_36) : $signed(_GEN_235); // @[CFARUtils.scala 433:24]
  assign _GEN_237 = 6'h25 == _T_8[5:0] ? $signed(adjShiftRegOut_37) : $signed(_GEN_236); // @[CFARUtils.scala 433:24]
  assign _GEN_238 = 6'h26 == _T_8[5:0] ? $signed(adjShiftRegOut_38) : $signed(_GEN_237); // @[CFARUtils.scala 433:24]
  assign _GEN_239 = 6'h27 == _T_8[5:0] ? $signed(adjShiftRegOut_39) : $signed(_GEN_238); // @[CFARUtils.scala 433:24]
  assign _GEN_240 = 6'h28 == _T_8[5:0] ? $signed(adjShiftRegOut_40) : $signed(_GEN_239); // @[CFARUtils.scala 433:24]
  assign _GEN_241 = 6'h29 == _T_8[5:0] ? $signed(adjShiftRegOut_41) : $signed(_GEN_240); // @[CFARUtils.scala 433:24]
  assign _GEN_242 = 6'h2a == _T_8[5:0] ? $signed(adjShiftRegOut_42) : $signed(_GEN_241); // @[CFARUtils.scala 433:24]
  assign _GEN_243 = 6'h2b == _T_8[5:0] ? $signed(adjShiftRegOut_43) : $signed(_GEN_242); // @[CFARUtils.scala 433:24]
  assign _GEN_244 = 6'h2c == _T_8[5:0] ? $signed(adjShiftRegOut_44) : $signed(_GEN_243); // @[CFARUtils.scala 433:24]
  assign _GEN_245 = 6'h2d == _T_8[5:0] ? $signed(adjShiftRegOut_45) : $signed(_GEN_244); // @[CFARUtils.scala 433:24]
  assign _GEN_246 = 6'h2e == _T_8[5:0] ? $signed(adjShiftRegOut_46) : $signed(_GEN_245); // @[CFARUtils.scala 433:24]
  assign _GEN_247 = 6'h2f == _T_8[5:0] ? $signed(adjShiftRegOut_47) : $signed(_GEN_246); // @[CFARUtils.scala 433:24]
  assign _GEN_248 = 6'h30 == _T_8[5:0] ? $signed(adjShiftRegOut_48) : $signed(_GEN_247); // @[CFARUtils.scala 433:24]
  assign _GEN_249 = 6'h31 == _T_8[5:0] ? $signed(adjShiftRegOut_49) : $signed(_GEN_248); // @[CFARUtils.scala 433:24]
  assign _GEN_250 = 6'h32 == _T_8[5:0] ? $signed(adjShiftRegOut_50) : $signed(_GEN_249); // @[CFARUtils.scala 433:24]
  assign _GEN_251 = 6'h33 == _T_8[5:0] ? $signed(adjShiftRegOut_51) : $signed(_GEN_250); // @[CFARUtils.scala 433:24]
  assign _GEN_252 = 6'h34 == _T_8[5:0] ? $signed(adjShiftRegOut_52) : $signed(_GEN_251); // @[CFARUtils.scala 433:24]
  assign _GEN_253 = 6'h35 == _T_8[5:0] ? $signed(adjShiftRegOut_53) : $signed(_GEN_252); // @[CFARUtils.scala 433:24]
  assign _GEN_254 = 6'h36 == _T_8[5:0] ? $signed(adjShiftRegOut_54) : $signed(_GEN_253); // @[CFARUtils.scala 433:24]
  assign _GEN_255 = 6'h37 == _T_8[5:0] ? $signed(adjShiftRegOut_55) : $signed(_GEN_254); // @[CFARUtils.scala 433:24]
  assign _GEN_256 = 6'h38 == _T_8[5:0] ? $signed(adjShiftRegOut_56) : $signed(_GEN_255); // @[CFARUtils.scala 433:24]
  assign _GEN_257 = 6'h39 == _T_8[5:0] ? $signed(adjShiftRegOut_57) : $signed(_GEN_256); // @[CFARUtils.scala 433:24]
  assign _GEN_258 = 6'h3a == _T_8[5:0] ? $signed(adjShiftRegOut_58) : $signed(_GEN_257); // @[CFARUtils.scala 433:24]
  assign _GEN_259 = 6'h3b == _T_8[5:0] ? $signed(adjShiftRegOut_59) : $signed(_GEN_258); // @[CFARUtils.scala 433:24]
  assign _GEN_260 = 6'h3c == _T_8[5:0] ? $signed(adjShiftRegOut_60) : $signed(_GEN_259); // @[CFARUtils.scala 433:24]
  assign _GEN_261 = 6'h3d == _T_8[5:0] ? $signed(adjShiftRegOut_61) : $signed(_GEN_260); // @[CFARUtils.scala 433:24]
  assign _GEN_262 = 6'h3e == _T_8[5:0] ? $signed(adjShiftRegOut_62) : $signed(_GEN_261); // @[CFARUtils.scala 433:24]
  assign _GEN_263 = 6'h3f == _T_8[5:0] ? $signed(adjShiftRegOut_63) : $signed(_GEN_262); // @[CFARUtils.scala 433:24]
  assign _T_823 = InitialInDone & io_in_valid; // @[CFARUtils.scala 436:70]
  assign _T_824 = last & en; // @[CFARUtils.scala 436:94]
  assign _T_825 = _T_823 | _T_824; // @[CFARUtils.scala 436:85]
  assign io_in_ready = _T_810 ? io_out_ready : _T_814; // @[CFARUtils.scala 426:20]
  assign io_out_valid = _T_810 ? io_in_valid : _T_825; // @[CFARUtils.scala 436:18]
  assign io_out_bits = _T_810 ? $signed(io_in_bits) : $signed(_GEN_263); // @[CFARUtils.scala 433:18]
  assign io_lastOut = _T_810 ? _T_395 : _GEN_196; // @[CFARUtils.scala 435:18]
  assign io_parallelOut_0 = adjShiftRegOut_0; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_1 = adjShiftRegOut_1; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_2 = adjShiftRegOut_2; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_3 = adjShiftRegOut_3; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_4 = adjShiftRegOut_4; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_5 = adjShiftRegOut_5; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_6 = adjShiftRegOut_6; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_7 = adjShiftRegOut_7; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_8 = adjShiftRegOut_8; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_9 = adjShiftRegOut_9; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_10 = adjShiftRegOut_10; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_11 = adjShiftRegOut_11; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_12 = adjShiftRegOut_12; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_13 = adjShiftRegOut_13; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_14 = adjShiftRegOut_14; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_15 = adjShiftRegOut_15; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_16 = adjShiftRegOut_16; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_17 = adjShiftRegOut_17; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_18 = adjShiftRegOut_18; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_19 = adjShiftRegOut_19; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_20 = adjShiftRegOut_20; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_21 = adjShiftRegOut_21; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_22 = adjShiftRegOut_22; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_23 = adjShiftRegOut_23; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_24 = adjShiftRegOut_24; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_25 = adjShiftRegOut_25; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_26 = adjShiftRegOut_26; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_27 = adjShiftRegOut_27; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_28 = adjShiftRegOut_28; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_29 = adjShiftRegOut_29; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_30 = adjShiftRegOut_30; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_31 = adjShiftRegOut_31; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_32 = adjShiftRegOut_32; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_33 = adjShiftRegOut_33; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_34 = adjShiftRegOut_34; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_35 = adjShiftRegOut_35; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_36 = adjShiftRegOut_36; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_37 = adjShiftRegOut_37; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_38 = adjShiftRegOut_38; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_39 = adjShiftRegOut_39; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_40 = adjShiftRegOut_40; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_41 = adjShiftRegOut_41; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_42 = adjShiftRegOut_42; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_43 = adjShiftRegOut_43; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_44 = adjShiftRegOut_44; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_45 = adjShiftRegOut_45; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_46 = adjShiftRegOut_46; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_47 = adjShiftRegOut_47; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_48 = adjShiftRegOut_48; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_49 = adjShiftRegOut_49; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_50 = adjShiftRegOut_50; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_51 = adjShiftRegOut_51; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_52 = adjShiftRegOut_52; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_53 = adjShiftRegOut_53; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_54 = adjShiftRegOut_54; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_55 = adjShiftRegOut_55; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_56 = adjShiftRegOut_56; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_57 = adjShiftRegOut_57; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_58 = adjShiftRegOut_58; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_59 = adjShiftRegOut_59; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_60 = adjShiftRegOut_60; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_61 = adjShiftRegOut_61; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_62 = adjShiftRegOut_62; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_63 = adjShiftRegOut_63; // @[CFARUtils.scala 434:18]
  assign io_cnt = cntIn; // @[CFARUtils.scala 438:16]
  assign io_regFull = InitialInDone & _T_808; // @[CFARUtils.scala 421:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  InitialInDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  last = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  adjShiftRegOut_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  adjShiftRegOut_1 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  adjShiftRegOut_2 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  adjShiftRegOut_3 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  adjShiftRegOut_4 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  adjShiftRegOut_5 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  adjShiftRegOut_6 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  adjShiftRegOut_7 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  adjShiftRegOut_8 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  adjShiftRegOut_9 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  adjShiftRegOut_10 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  adjShiftRegOut_11 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  adjShiftRegOut_12 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  adjShiftRegOut_13 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  adjShiftRegOut_14 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  adjShiftRegOut_15 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  adjShiftRegOut_16 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  adjShiftRegOut_17 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  adjShiftRegOut_18 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  adjShiftRegOut_19 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  adjShiftRegOut_20 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  adjShiftRegOut_21 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  adjShiftRegOut_22 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  adjShiftRegOut_23 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  adjShiftRegOut_24 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  adjShiftRegOut_25 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  adjShiftRegOut_26 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  adjShiftRegOut_27 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  adjShiftRegOut_28 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  adjShiftRegOut_29 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  adjShiftRegOut_30 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  adjShiftRegOut_31 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  adjShiftRegOut_32 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  adjShiftRegOut_33 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  adjShiftRegOut_34 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  adjShiftRegOut_35 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  adjShiftRegOut_36 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  adjShiftRegOut_37 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  adjShiftRegOut_38 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  adjShiftRegOut_39 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  adjShiftRegOut_40 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  adjShiftRegOut_41 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  adjShiftRegOut_42 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  adjShiftRegOut_43 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  adjShiftRegOut_44 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  adjShiftRegOut_45 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  adjShiftRegOut_46 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  adjShiftRegOut_47 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  adjShiftRegOut_48 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  adjShiftRegOut_49 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  adjShiftRegOut_50 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  adjShiftRegOut_51 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  adjShiftRegOut_52 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  adjShiftRegOut_53 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  adjShiftRegOut_54 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  adjShiftRegOut_55 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  adjShiftRegOut_56 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  adjShiftRegOut_57 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  adjShiftRegOut_58 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  adjShiftRegOut_59 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  adjShiftRegOut_60 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  adjShiftRegOut_61 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  adjShiftRegOut_62 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  adjShiftRegOut_63 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  cntIn = _RAND_66[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_736 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_737 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_738 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_739 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_740 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_741 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_742 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_743 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_744 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_745 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_746 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_747 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_748 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_749 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_750 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_751 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_752 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_753 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_754 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_755 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_756 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_757 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_758 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_759 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_760 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_761 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_762 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_763 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_764 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_765 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_766 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_767 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_768 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_769 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_770 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_771 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_772 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_773 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_774 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_775 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_776 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_777 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_778 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_779 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_780 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_781 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_782 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_783 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_784 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_785 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_786 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_787 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_788 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_789 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_790 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_791 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_792 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_793 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_794 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_795 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_796 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_797 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_798 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_799 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      InitialInDone <= 1'h0;
    end else if (_T_804) begin
      InitialInDone <= 1'h0;
    end else if (_T_399) begin
      InitialInDone <= _GEN_66;
    end else begin
      InitialInDone <= _GEN_67;
    end
    if (reset) begin
      last <= 1'h0;
    end else if (_T_804) begin
      last <= 1'h0;
    end else begin
      last <= _GEN_64;
    end
    if (reset) begin
      adjShiftRegOut_0 <= 16'sh0;
    end else if (_T_326) begin
      adjShiftRegOut_0 <= io_in_bits;
    end
    if (reset) begin
      adjShiftRegOut_1 <= 16'sh0;
    end else if (_T_325) begin
      adjShiftRegOut_1 <= adjShiftRegOut_0;
    end
    if (reset) begin
      adjShiftRegOut_2 <= 16'sh0;
    end else if (_T_324) begin
      adjShiftRegOut_2 <= adjShiftRegOut_1;
    end
    if (reset) begin
      adjShiftRegOut_3 <= 16'sh0;
    end else if (_T_323) begin
      adjShiftRegOut_3 <= adjShiftRegOut_2;
    end
    if (reset) begin
      adjShiftRegOut_4 <= 16'sh0;
    end else if (_T_322) begin
      adjShiftRegOut_4 <= adjShiftRegOut_3;
    end
    if (reset) begin
      adjShiftRegOut_5 <= 16'sh0;
    end else if (_T_321) begin
      adjShiftRegOut_5 <= adjShiftRegOut_4;
    end
    if (reset) begin
      adjShiftRegOut_6 <= 16'sh0;
    end else if (_T_320) begin
      adjShiftRegOut_6 <= adjShiftRegOut_5;
    end
    if (reset) begin
      adjShiftRegOut_7 <= 16'sh0;
    end else if (_T_319) begin
      adjShiftRegOut_7 <= adjShiftRegOut_6;
    end
    if (reset) begin
      adjShiftRegOut_8 <= 16'sh0;
    end else if (_T_318) begin
      adjShiftRegOut_8 <= adjShiftRegOut_7;
    end
    if (reset) begin
      adjShiftRegOut_9 <= 16'sh0;
    end else if (_T_317) begin
      adjShiftRegOut_9 <= adjShiftRegOut_8;
    end
    if (reset) begin
      adjShiftRegOut_10 <= 16'sh0;
    end else if (_T_316) begin
      adjShiftRegOut_10 <= adjShiftRegOut_9;
    end
    if (reset) begin
      adjShiftRegOut_11 <= 16'sh0;
    end else if (_T_315) begin
      adjShiftRegOut_11 <= adjShiftRegOut_10;
    end
    if (reset) begin
      adjShiftRegOut_12 <= 16'sh0;
    end else if (_T_314) begin
      adjShiftRegOut_12 <= adjShiftRegOut_11;
    end
    if (reset) begin
      adjShiftRegOut_13 <= 16'sh0;
    end else if (_T_313) begin
      adjShiftRegOut_13 <= adjShiftRegOut_12;
    end
    if (reset) begin
      adjShiftRegOut_14 <= 16'sh0;
    end else if (_T_312) begin
      adjShiftRegOut_14 <= adjShiftRegOut_13;
    end
    if (reset) begin
      adjShiftRegOut_15 <= 16'sh0;
    end else if (_T_311) begin
      adjShiftRegOut_15 <= adjShiftRegOut_14;
    end
    if (reset) begin
      adjShiftRegOut_16 <= 16'sh0;
    end else if (_T_310) begin
      adjShiftRegOut_16 <= adjShiftRegOut_15;
    end
    if (reset) begin
      adjShiftRegOut_17 <= 16'sh0;
    end else if (_T_309) begin
      adjShiftRegOut_17 <= adjShiftRegOut_16;
    end
    if (reset) begin
      adjShiftRegOut_18 <= 16'sh0;
    end else if (_T_308) begin
      adjShiftRegOut_18 <= adjShiftRegOut_17;
    end
    if (reset) begin
      adjShiftRegOut_19 <= 16'sh0;
    end else if (_T_307) begin
      adjShiftRegOut_19 <= adjShiftRegOut_18;
    end
    if (reset) begin
      adjShiftRegOut_20 <= 16'sh0;
    end else if (_T_306) begin
      adjShiftRegOut_20 <= adjShiftRegOut_19;
    end
    if (reset) begin
      adjShiftRegOut_21 <= 16'sh0;
    end else if (_T_305) begin
      adjShiftRegOut_21 <= adjShiftRegOut_20;
    end
    if (reset) begin
      adjShiftRegOut_22 <= 16'sh0;
    end else if (_T_304) begin
      adjShiftRegOut_22 <= adjShiftRegOut_21;
    end
    if (reset) begin
      adjShiftRegOut_23 <= 16'sh0;
    end else if (_T_303) begin
      adjShiftRegOut_23 <= adjShiftRegOut_22;
    end
    if (reset) begin
      adjShiftRegOut_24 <= 16'sh0;
    end else if (_T_302) begin
      adjShiftRegOut_24 <= adjShiftRegOut_23;
    end
    if (reset) begin
      adjShiftRegOut_25 <= 16'sh0;
    end else if (_T_301) begin
      adjShiftRegOut_25 <= adjShiftRegOut_24;
    end
    if (reset) begin
      adjShiftRegOut_26 <= 16'sh0;
    end else if (_T_300) begin
      adjShiftRegOut_26 <= adjShiftRegOut_25;
    end
    if (reset) begin
      adjShiftRegOut_27 <= 16'sh0;
    end else if (_T_299) begin
      adjShiftRegOut_27 <= adjShiftRegOut_26;
    end
    if (reset) begin
      adjShiftRegOut_28 <= 16'sh0;
    end else if (_T_298) begin
      adjShiftRegOut_28 <= adjShiftRegOut_27;
    end
    if (reset) begin
      adjShiftRegOut_29 <= 16'sh0;
    end else if (_T_297) begin
      adjShiftRegOut_29 <= adjShiftRegOut_28;
    end
    if (reset) begin
      adjShiftRegOut_30 <= 16'sh0;
    end else if (_T_296) begin
      adjShiftRegOut_30 <= adjShiftRegOut_29;
    end
    if (reset) begin
      adjShiftRegOut_31 <= 16'sh0;
    end else if (_T_295) begin
      adjShiftRegOut_31 <= adjShiftRegOut_30;
    end
    if (reset) begin
      adjShiftRegOut_32 <= 16'sh0;
    end else if (_T_294) begin
      adjShiftRegOut_32 <= adjShiftRegOut_31;
    end
    if (reset) begin
      adjShiftRegOut_33 <= 16'sh0;
    end else if (_T_293) begin
      adjShiftRegOut_33 <= adjShiftRegOut_32;
    end
    if (reset) begin
      adjShiftRegOut_34 <= 16'sh0;
    end else if (_T_292) begin
      adjShiftRegOut_34 <= adjShiftRegOut_33;
    end
    if (reset) begin
      adjShiftRegOut_35 <= 16'sh0;
    end else if (_T_291) begin
      adjShiftRegOut_35 <= adjShiftRegOut_34;
    end
    if (reset) begin
      adjShiftRegOut_36 <= 16'sh0;
    end else if (_T_290) begin
      adjShiftRegOut_36 <= adjShiftRegOut_35;
    end
    if (reset) begin
      adjShiftRegOut_37 <= 16'sh0;
    end else if (_T_289) begin
      adjShiftRegOut_37 <= adjShiftRegOut_36;
    end
    if (reset) begin
      adjShiftRegOut_38 <= 16'sh0;
    end else if (_T_288) begin
      adjShiftRegOut_38 <= adjShiftRegOut_37;
    end
    if (reset) begin
      adjShiftRegOut_39 <= 16'sh0;
    end else if (_T_287) begin
      adjShiftRegOut_39 <= adjShiftRegOut_38;
    end
    if (reset) begin
      adjShiftRegOut_40 <= 16'sh0;
    end else if (_T_286) begin
      adjShiftRegOut_40 <= adjShiftRegOut_39;
    end
    if (reset) begin
      adjShiftRegOut_41 <= 16'sh0;
    end else if (_T_285) begin
      adjShiftRegOut_41 <= adjShiftRegOut_40;
    end
    if (reset) begin
      adjShiftRegOut_42 <= 16'sh0;
    end else if (_T_284) begin
      adjShiftRegOut_42 <= adjShiftRegOut_41;
    end
    if (reset) begin
      adjShiftRegOut_43 <= 16'sh0;
    end else if (_T_283) begin
      adjShiftRegOut_43 <= adjShiftRegOut_42;
    end
    if (reset) begin
      adjShiftRegOut_44 <= 16'sh0;
    end else if (_T_282) begin
      adjShiftRegOut_44 <= adjShiftRegOut_43;
    end
    if (reset) begin
      adjShiftRegOut_45 <= 16'sh0;
    end else if (_T_281) begin
      adjShiftRegOut_45 <= adjShiftRegOut_44;
    end
    if (reset) begin
      adjShiftRegOut_46 <= 16'sh0;
    end else if (_T_280) begin
      adjShiftRegOut_46 <= adjShiftRegOut_45;
    end
    if (reset) begin
      adjShiftRegOut_47 <= 16'sh0;
    end else if (_T_279) begin
      adjShiftRegOut_47 <= adjShiftRegOut_46;
    end
    if (reset) begin
      adjShiftRegOut_48 <= 16'sh0;
    end else if (_T_278) begin
      adjShiftRegOut_48 <= adjShiftRegOut_47;
    end
    if (reset) begin
      adjShiftRegOut_49 <= 16'sh0;
    end else if (_T_277) begin
      adjShiftRegOut_49 <= adjShiftRegOut_48;
    end
    if (reset) begin
      adjShiftRegOut_50 <= 16'sh0;
    end else if (_T_276) begin
      adjShiftRegOut_50 <= adjShiftRegOut_49;
    end
    if (reset) begin
      adjShiftRegOut_51 <= 16'sh0;
    end else if (_T_275) begin
      adjShiftRegOut_51 <= adjShiftRegOut_50;
    end
    if (reset) begin
      adjShiftRegOut_52 <= 16'sh0;
    end else if (_T_274) begin
      adjShiftRegOut_52 <= adjShiftRegOut_51;
    end
    if (reset) begin
      adjShiftRegOut_53 <= 16'sh0;
    end else if (_T_273) begin
      adjShiftRegOut_53 <= adjShiftRegOut_52;
    end
    if (reset) begin
      adjShiftRegOut_54 <= 16'sh0;
    end else if (_T_272) begin
      adjShiftRegOut_54 <= adjShiftRegOut_53;
    end
    if (reset) begin
      adjShiftRegOut_55 <= 16'sh0;
    end else if (_T_271) begin
      adjShiftRegOut_55 <= adjShiftRegOut_54;
    end
    if (reset) begin
      adjShiftRegOut_56 <= 16'sh0;
    end else if (_T_270) begin
      adjShiftRegOut_56 <= adjShiftRegOut_55;
    end
    if (reset) begin
      adjShiftRegOut_57 <= 16'sh0;
    end else if (_T_269) begin
      adjShiftRegOut_57 <= adjShiftRegOut_56;
    end
    if (reset) begin
      adjShiftRegOut_58 <= 16'sh0;
    end else if (_T_268) begin
      adjShiftRegOut_58 <= adjShiftRegOut_57;
    end
    if (reset) begin
      adjShiftRegOut_59 <= 16'sh0;
    end else if (_T_267) begin
      adjShiftRegOut_59 <= adjShiftRegOut_58;
    end
    if (reset) begin
      adjShiftRegOut_60 <= 16'sh0;
    end else if (_T_266) begin
      adjShiftRegOut_60 <= adjShiftRegOut_59;
    end
    if (reset) begin
      adjShiftRegOut_61 <= 16'sh0;
    end else if (_T_265) begin
      adjShiftRegOut_61 <= adjShiftRegOut_60;
    end
    if (reset) begin
      adjShiftRegOut_62 <= 16'sh0;
    end else if (_T_264) begin
      adjShiftRegOut_62 <= adjShiftRegOut_61;
    end
    if (reset) begin
      adjShiftRegOut_63 <= 16'sh0;
    end else if (_T_263) begin
      adjShiftRegOut_63 <= adjShiftRegOut_62;
    end
    if (reset) begin
      cntIn <= 7'h0;
    end else if (_T_804) begin
      cntIn <= 7'h0;
    end else if (_T_1) begin
      cntIn <= _T_398;
    end
    if (reset) begin
      _T_736 <= 1'h0;
    end else if (_T_409) begin
      _T_736 <= _T_395;
    end
    if (reset) begin
      _T_737 <= 1'h0;
    end else if (_T_734) begin
      _T_737 <= _T_736;
    end
    if (reset) begin
      _T_738 <= 1'h0;
    end else if (_T_733) begin
      _T_738 <= _T_737;
    end
    if (reset) begin
      _T_739 <= 1'h0;
    end else if (_T_732) begin
      _T_739 <= _T_738;
    end
    if (reset) begin
      _T_740 <= 1'h0;
    end else if (_T_731) begin
      _T_740 <= _T_739;
    end
    if (reset) begin
      _T_741 <= 1'h0;
    end else if (_T_730) begin
      _T_741 <= _T_740;
    end
    if (reset) begin
      _T_742 <= 1'h0;
    end else if (_T_729) begin
      _T_742 <= _T_741;
    end
    if (reset) begin
      _T_743 <= 1'h0;
    end else if (_T_728) begin
      _T_743 <= _T_742;
    end
    if (reset) begin
      _T_744 <= 1'h0;
    end else if (_T_727) begin
      _T_744 <= _T_743;
    end
    if (reset) begin
      _T_745 <= 1'h0;
    end else if (_T_726) begin
      _T_745 <= _T_744;
    end
    if (reset) begin
      _T_746 <= 1'h0;
    end else if (_T_725) begin
      _T_746 <= _T_745;
    end
    if (reset) begin
      _T_747 <= 1'h0;
    end else if (_T_724) begin
      _T_747 <= _T_746;
    end
    if (reset) begin
      _T_748 <= 1'h0;
    end else if (_T_723) begin
      _T_748 <= _T_747;
    end
    if (reset) begin
      _T_749 <= 1'h0;
    end else if (_T_722) begin
      _T_749 <= _T_748;
    end
    if (reset) begin
      _T_750 <= 1'h0;
    end else if (_T_721) begin
      _T_750 <= _T_749;
    end
    if (reset) begin
      _T_751 <= 1'h0;
    end else if (_T_720) begin
      _T_751 <= _T_750;
    end
    if (reset) begin
      _T_752 <= 1'h0;
    end else if (_T_719) begin
      _T_752 <= _T_751;
    end
    if (reset) begin
      _T_753 <= 1'h0;
    end else if (_T_718) begin
      _T_753 <= _T_752;
    end
    if (reset) begin
      _T_754 <= 1'h0;
    end else if (_T_717) begin
      _T_754 <= _T_753;
    end
    if (reset) begin
      _T_755 <= 1'h0;
    end else if (_T_716) begin
      _T_755 <= _T_754;
    end
    if (reset) begin
      _T_756 <= 1'h0;
    end else if (_T_715) begin
      _T_756 <= _T_755;
    end
    if (reset) begin
      _T_757 <= 1'h0;
    end else if (_T_714) begin
      _T_757 <= _T_756;
    end
    if (reset) begin
      _T_758 <= 1'h0;
    end else if (_T_713) begin
      _T_758 <= _T_757;
    end
    if (reset) begin
      _T_759 <= 1'h0;
    end else if (_T_712) begin
      _T_759 <= _T_758;
    end
    if (reset) begin
      _T_760 <= 1'h0;
    end else if (_T_711) begin
      _T_760 <= _T_759;
    end
    if (reset) begin
      _T_761 <= 1'h0;
    end else if (_T_710) begin
      _T_761 <= _T_760;
    end
    if (reset) begin
      _T_762 <= 1'h0;
    end else if (_T_709) begin
      _T_762 <= _T_761;
    end
    if (reset) begin
      _T_763 <= 1'h0;
    end else if (_T_708) begin
      _T_763 <= _T_762;
    end
    if (reset) begin
      _T_764 <= 1'h0;
    end else if (_T_707) begin
      _T_764 <= _T_763;
    end
    if (reset) begin
      _T_765 <= 1'h0;
    end else if (_T_706) begin
      _T_765 <= _T_764;
    end
    if (reset) begin
      _T_766 <= 1'h0;
    end else if (_T_705) begin
      _T_766 <= _T_765;
    end
    if (reset) begin
      _T_767 <= 1'h0;
    end else if (_T_704) begin
      _T_767 <= _T_766;
    end
    if (reset) begin
      _T_768 <= 1'h0;
    end else if (_T_703) begin
      _T_768 <= _T_767;
    end
    if (reset) begin
      _T_769 <= 1'h0;
    end else if (_T_702) begin
      _T_769 <= _T_768;
    end
    if (reset) begin
      _T_770 <= 1'h0;
    end else if (_T_701) begin
      _T_770 <= _T_769;
    end
    if (reset) begin
      _T_771 <= 1'h0;
    end else if (_T_700) begin
      _T_771 <= _T_770;
    end
    if (reset) begin
      _T_772 <= 1'h0;
    end else if (_T_699) begin
      _T_772 <= _T_771;
    end
    if (reset) begin
      _T_773 <= 1'h0;
    end else if (_T_698) begin
      _T_773 <= _T_772;
    end
    if (reset) begin
      _T_774 <= 1'h0;
    end else if (_T_697) begin
      _T_774 <= _T_773;
    end
    if (reset) begin
      _T_775 <= 1'h0;
    end else if (_T_696) begin
      _T_775 <= _T_774;
    end
    if (reset) begin
      _T_776 <= 1'h0;
    end else if (_T_695) begin
      _T_776 <= _T_775;
    end
    if (reset) begin
      _T_777 <= 1'h0;
    end else if (_T_694) begin
      _T_777 <= _T_776;
    end
    if (reset) begin
      _T_778 <= 1'h0;
    end else if (_T_693) begin
      _T_778 <= _T_777;
    end
    if (reset) begin
      _T_779 <= 1'h0;
    end else if (_T_692) begin
      _T_779 <= _T_778;
    end
    if (reset) begin
      _T_780 <= 1'h0;
    end else if (_T_691) begin
      _T_780 <= _T_779;
    end
    if (reset) begin
      _T_781 <= 1'h0;
    end else if (_T_690) begin
      _T_781 <= _T_780;
    end
    if (reset) begin
      _T_782 <= 1'h0;
    end else if (_T_689) begin
      _T_782 <= _T_781;
    end
    if (reset) begin
      _T_783 <= 1'h0;
    end else if (_T_688) begin
      _T_783 <= _T_782;
    end
    if (reset) begin
      _T_784 <= 1'h0;
    end else if (_T_687) begin
      _T_784 <= _T_783;
    end
    if (reset) begin
      _T_785 <= 1'h0;
    end else if (_T_686) begin
      _T_785 <= _T_784;
    end
    if (reset) begin
      _T_786 <= 1'h0;
    end else if (_T_685) begin
      _T_786 <= _T_785;
    end
    if (reset) begin
      _T_787 <= 1'h0;
    end else if (_T_684) begin
      _T_787 <= _T_786;
    end
    if (reset) begin
      _T_788 <= 1'h0;
    end else if (_T_683) begin
      _T_788 <= _T_787;
    end
    if (reset) begin
      _T_789 <= 1'h0;
    end else if (_T_682) begin
      _T_789 <= _T_788;
    end
    if (reset) begin
      _T_790 <= 1'h0;
    end else if (_T_681) begin
      _T_790 <= _T_789;
    end
    if (reset) begin
      _T_791 <= 1'h0;
    end else if (_T_680) begin
      _T_791 <= _T_790;
    end
    if (reset) begin
      _T_792 <= 1'h0;
    end else if (_T_679) begin
      _T_792 <= _T_791;
    end
    if (reset) begin
      _T_793 <= 1'h0;
    end else if (_T_678) begin
      _T_793 <= _T_792;
    end
    if (reset) begin
      _T_794 <= 1'h0;
    end else if (_T_677) begin
      _T_794 <= _T_793;
    end
    if (reset) begin
      _T_795 <= 1'h0;
    end else if (_T_676) begin
      _T_795 <= _T_794;
    end
    if (reset) begin
      _T_796 <= 1'h0;
    end else if (_T_675) begin
      _T_796 <= _T_795;
    end
    if (reset) begin
      _T_797 <= 1'h0;
    end else if (_T_674) begin
      _T_797 <= _T_796;
    end
    if (reset) begin
      _T_798 <= 1'h0;
    end else if (_T_673) begin
      _T_798 <= _T_797;
    end
    if (reset) begin
      _T_799 <= 1'h0;
    end else if (_T_672) begin
      _T_799 <= _T_798;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:345 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 345:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[CFARUtils.scala 345:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:330 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 330:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[CFARUtils.scala 330:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AdjustableShiftRegisterStream_1(
  input         clock,
  input         reset,
  input  [3:0]  io_depth,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut,
  output [15:0] io_parallelOut_0,
  output [15:0] io_parallelOut_1,
  output [15:0] io_parallelOut_2,
  output [15:0] io_parallelOut_3,
  output [15:0] io_parallelOut_4,
  output [15:0] io_parallelOut_5,
  output [15:0] io_parallelOut_6,
  output [15:0] io_parallelOut_7
);
  reg  InitialInDone; // @[CFARUtils.scala 379:30]
  reg [31:0] _RAND_0;
  reg  last; // @[CFARUtils.scala 380:21]
  reg [31:0] _RAND_1;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[CFARUtils.scala 385:34]
  wire  en; // @[CFARUtils.scala 385:25]
  wire  _T_3; // @[CFARUtils.scala 345:18]
  wire  _T_5; // @[CFARUtils.scala 345:11]
  wire  _T_6; // @[CFARUtils.scala 345:11]
  wire [3:0] _T_8; // @[CFARUtils.scala 350:87]
  wire  _T_9; // @[CFARUtils.scala 350:78]
  wire  _T_13; // @[CFARUtils.scala 350:78]
  wire  _T_14; // @[CFARUtils.scala 350:94]
  wire  _T_17; // @[CFARUtils.scala 350:78]
  wire  _T_18; // @[CFARUtils.scala 350:94]
  wire  _T_21; // @[CFARUtils.scala 350:78]
  wire  _T_22; // @[CFARUtils.scala 350:94]
  wire  _T_25; // @[CFARUtils.scala 350:78]
  wire  _T_26; // @[CFARUtils.scala 350:94]
  wire  _T_29; // @[CFARUtils.scala 350:78]
  wire  _T_30; // @[CFARUtils.scala 350:94]
  wire  _T_33; // @[CFARUtils.scala 350:78]
  wire  _T_34; // @[CFARUtils.scala 350:94]
  wire  _T_37; // @[CFARUtils.scala 350:78]
  wire  _T_38; // @[CFARUtils.scala 350:94]
  wire  activeRegs_7; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_39; // @[CFARUtils.scala 319:37]
  wire  activeRegs_6; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_40; // @[CFARUtils.scala 319:37]
  wire  activeRegs_5; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_41; // @[CFARUtils.scala 319:37]
  wire  activeRegs_4; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_42; // @[CFARUtils.scala 319:37]
  wire  activeRegs_3; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_43; // @[CFARUtils.scala 319:37]
  wire  activeRegs_2; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_44; // @[CFARUtils.scala 319:37]
  wire  activeRegs_1; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_45; // @[CFARUtils.scala 319:37]
  wire  activeRegs_0; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_46; // @[CFARUtils.scala 319:37]
  reg [15:0] adjShiftRegOut_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [15:0] adjShiftRegOut_1; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [15:0] adjShiftRegOut_2; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [15:0] adjShiftRegOut_3; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [15:0] adjShiftRegOut_4; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [15:0] adjShiftRegOut_5; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [15:0] adjShiftRegOut_6; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  reg [15:0] adjShiftRegOut_7; // @[Reg.scala 27:20]
  reg [31:0] _RAND_9;
  reg [3:0] cntIn; // @[CFARUtils.scala 390:23]
  reg [31:0] _RAND_10;
  wire  _T_59; // @[CFARUtils.scala 392:19]
  wire  _GEN_8; // @[CFARUtils.scala 392:36]
  wire [3:0] _T_62; // @[CFARUtils.scala 397:20]
  wire  _T_63; // @[CFARUtils.scala 400:18]
  wire  _T_66; // @[CFARUtils.scala 401:17]
  wire  _T_68; // @[CFARUtils.scala 401:36]
  wire  _GEN_10; // @[CFARUtils.scala 401:53]
  wire  _T_70; // @[CFARUtils.scala 406:36]
  wire  _T_71; // @[CFARUtils.scala 406:24]
  wire  _GEN_11; // @[CFARUtils.scala 406:45]
  wire  _T_73; // @[Decoupled.scala 40:37]
  wire  _T_112; // @[CFARUtils.scala 319:37]
  wire  _T_113; // @[CFARUtils.scala 319:37]
  wire  _T_114; // @[CFARUtils.scala 319:37]
  wire  _T_115; // @[CFARUtils.scala 319:37]
  wire  _T_116; // @[CFARUtils.scala 319:37]
  wire  _T_117; // @[CFARUtils.scala 319:37]
  wire  _T_118; // @[CFARUtils.scala 319:37]
  reg  _T_120; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg  _T_121; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg  _T_122; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg  _T_123; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  reg  _T_124; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  reg  _T_125; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg  _T_126; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  reg  _T_127; // @[Reg.scala 27:20]
  reg [31:0] _RAND_18;
  wire  _GEN_22; // @[CFARUtils.scala 414:17]
  wire  _GEN_23; // @[CFARUtils.scala 414:17]
  wire  _GEN_24; // @[CFARUtils.scala 414:17]
  wire  _GEN_25; // @[CFARUtils.scala 414:17]
  wire  _GEN_26; // @[CFARUtils.scala 414:17]
  wire  _GEN_27; // @[CFARUtils.scala 414:17]
  wire  _GEN_28; // @[CFARUtils.scala 414:17]
  wire  _T_132; // @[CFARUtils.scala 414:17]
  wire  _T_134; // @[CFARUtils.scala 420:36]
  wire  _T_136; // @[CFARUtils.scala 421:36]
  wire  _T_138; // @[CFARUtils.scala 426:37]
  wire  _T_141; // @[CFARUtils.scala 426:91]
  wire  _T_142; // @[CFARUtils.scala 426:75]
  wire [15:0] _GEN_33; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_34; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_35; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_36; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_37; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_38; // @[CFARUtils.scala 433:24]
  wire [15:0] _GEN_39; // @[CFARUtils.scala 433:24]
  wire  _T_151; // @[CFARUtils.scala 436:70]
  wire  _T_152; // @[CFARUtils.scala 436:94]
  wire  _T_153; // @[CFARUtils.scala 436:85]
  assign _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = last & io_out_ready; // @[CFARUtils.scala 385:34]
  assign en = _T_1 | _T_2; // @[CFARUtils.scala 385:25]
  assign _T_3 = io_depth <= 4'h8; // @[CFARUtils.scala 345:18]
  assign _T_5 = _T_3 | reset; // @[CFARUtils.scala 345:11]
  assign _T_6 = ~_T_5; // @[CFARUtils.scala 345:11]
  assign _T_8 = io_depth - 4'h1; // @[CFARUtils.scala 350:87]
  assign _T_9 = 1'h1; // @[CFARUtils.scala 350:78]
  assign _T_13 = 4'h1 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_14 = _T_13; // @[CFARUtils.scala 350:94]
  assign _T_17 = 4'h2 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_18 = _T_17; // @[CFARUtils.scala 350:94]
  assign _T_21 = 4'h3 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_22 = _T_21; // @[CFARUtils.scala 350:94]
  assign _T_25 = 4'h4 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_26 = _T_25; // @[CFARUtils.scala 350:94]
  assign _T_29 = 4'h5 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_30 = _T_29; // @[CFARUtils.scala 350:94]
  assign _T_33 = 4'h6 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_34 = _T_33; // @[CFARUtils.scala 350:94]
  assign _T_37 = 4'h7 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_38 = _T_37; // @[CFARUtils.scala 350:94]
  assign activeRegs_7 = _T_37; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_39 = _T_38 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_6 = _T_33; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_40 = _T_34 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_5 = _T_29; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_41 = _T_30 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_4 = _T_25; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_42 = _T_26 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_3 = _T_21; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_43 = _T_22 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_2 = _T_17; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_44 = _T_18 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_1 = _T_13; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_45 = _T_14 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_0 = 1'h1; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_46 = _T_9 & en; // @[CFARUtils.scala 319:37]
  assign _T_59 = io_lastIn & _T_1; // @[CFARUtils.scala 392:19]
  assign _GEN_8 = _T_59 | last; // @[CFARUtils.scala 392:36]
  assign _T_62 = cntIn + 4'h1; // @[CFARUtils.scala 397:20]
  assign _T_63 = io_depth > 4'h1; // @[CFARUtils.scala 400:18]
  assign _T_66 = cntIn == _T_8; // @[CFARUtils.scala 401:17]
  assign _T_68 = _T_66 & _T_1; // @[CFARUtils.scala 401:36]
  assign _GEN_10 = _T_68 | InitialInDone; // @[CFARUtils.scala 401:53]
  assign _T_70 = io_depth == 4'h1; // @[CFARUtils.scala 406:36]
  assign _T_71 = _T_1 & _T_70; // @[CFARUtils.scala 406:24]
  assign _GEN_11 = _T_71 | InitialInDone; // @[CFARUtils.scala 406:45]
  assign _T_73 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_112 = _T_37 & _T_73; // @[CFARUtils.scala 319:37]
  assign _T_113 = _T_33 & _T_73; // @[CFARUtils.scala 319:37]
  assign _T_114 = _T_29 & _T_73; // @[CFARUtils.scala 319:37]
  assign _T_115 = _T_25 & _T_73; // @[CFARUtils.scala 319:37]
  assign _T_116 = _T_21 & _T_73; // @[CFARUtils.scala 319:37]
  assign _T_117 = _T_17 & _T_73; // @[CFARUtils.scala 319:37]
  assign _T_118 = _T_13 & _T_73; // @[CFARUtils.scala 319:37]
  assign _GEN_22 = 3'h1 == _T_8[2:0] ? _T_121 : _T_120; // @[CFARUtils.scala 414:17]
  assign _GEN_23 = 3'h2 == _T_8[2:0] ? _T_122 : _GEN_22; // @[CFARUtils.scala 414:17]
  assign _GEN_24 = 3'h3 == _T_8[2:0] ? _T_123 : _GEN_23; // @[CFARUtils.scala 414:17]
  assign _GEN_25 = 3'h4 == _T_8[2:0] ? _T_124 : _GEN_24; // @[CFARUtils.scala 414:17]
  assign _GEN_26 = 3'h5 == _T_8[2:0] ? _T_125 : _GEN_25; // @[CFARUtils.scala 414:17]
  assign _GEN_27 = 3'h6 == _T_8[2:0] ? _T_126 : _GEN_26; // @[CFARUtils.scala 414:17]
  assign _GEN_28 = 3'h7 == _T_8[2:0] ? _T_127 : _GEN_27; // @[CFARUtils.scala 414:17]
  assign _T_132 = _GEN_28 & _T_73; // @[CFARUtils.scala 414:17]
  assign _T_134 = ~InitialInDone; // @[CFARUtils.scala 420:36]
  assign _T_136 = ~last; // @[CFARUtils.scala 421:36]
  assign _T_138 = io_depth == 4'h0; // @[CFARUtils.scala 426:37]
  assign _T_141 = io_out_ready & _T_136; // @[CFARUtils.scala 426:91]
  assign _T_142 = _T_134 | _T_141; // @[CFARUtils.scala 426:75]
  assign _GEN_33 = 3'h1 == _T_8[2:0] ? $signed(adjShiftRegOut_1) : $signed(adjShiftRegOut_0); // @[CFARUtils.scala 433:24]
  assign _GEN_34 = 3'h2 == _T_8[2:0] ? $signed(adjShiftRegOut_2) : $signed(_GEN_33); // @[CFARUtils.scala 433:24]
  assign _GEN_35 = 3'h3 == _T_8[2:0] ? $signed(adjShiftRegOut_3) : $signed(_GEN_34); // @[CFARUtils.scala 433:24]
  assign _GEN_36 = 3'h4 == _T_8[2:0] ? $signed(adjShiftRegOut_4) : $signed(_GEN_35); // @[CFARUtils.scala 433:24]
  assign _GEN_37 = 3'h5 == _T_8[2:0] ? $signed(adjShiftRegOut_5) : $signed(_GEN_36); // @[CFARUtils.scala 433:24]
  assign _GEN_38 = 3'h6 == _T_8[2:0] ? $signed(adjShiftRegOut_6) : $signed(_GEN_37); // @[CFARUtils.scala 433:24]
  assign _GEN_39 = 3'h7 == _T_8[2:0] ? $signed(adjShiftRegOut_7) : $signed(_GEN_38); // @[CFARUtils.scala 433:24]
  assign _T_151 = InitialInDone & io_in_valid; // @[CFARUtils.scala 436:70]
  assign _T_152 = last & en; // @[CFARUtils.scala 436:94]
  assign _T_153 = _T_151 | _T_152; // @[CFARUtils.scala 436:85]
  assign io_in_ready = _T_138 ? io_out_ready : _T_142; // @[CFARUtils.scala 426:20]
  assign io_out_valid = _T_138 ? io_in_valid : _T_153; // @[CFARUtils.scala 436:18]
  assign io_out_bits = _T_138 ? $signed(io_in_bits) : $signed(_GEN_39); // @[CFARUtils.scala 433:18]
  assign io_lastOut = _T_138 ? _T_59 : _GEN_28; // @[CFARUtils.scala 435:18]
  assign io_parallelOut_0 = adjShiftRegOut_0; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_1 = adjShiftRegOut_1; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_2 = adjShiftRegOut_2; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_3 = adjShiftRegOut_3; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_4 = adjShiftRegOut_4; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_5 = adjShiftRegOut_5; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_6 = adjShiftRegOut_6; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_7 = adjShiftRegOut_7; // @[CFARUtils.scala 434:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  InitialInDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  last = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  adjShiftRegOut_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  adjShiftRegOut_1 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  adjShiftRegOut_2 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  adjShiftRegOut_3 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  adjShiftRegOut_4 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  adjShiftRegOut_5 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  adjShiftRegOut_6 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  adjShiftRegOut_7 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  cntIn = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_120 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_121 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_122 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_123 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_124 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_125 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_126 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_127 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      InitialInDone <= 1'h0;
    end else if (_T_132) begin
      InitialInDone <= 1'h0;
    end else if (_T_63) begin
      InitialInDone <= _GEN_10;
    end else begin
      InitialInDone <= _GEN_11;
    end
    if (reset) begin
      last <= 1'h0;
    end else if (_T_132) begin
      last <= 1'h0;
    end else begin
      last <= _GEN_8;
    end
    if (reset) begin
      adjShiftRegOut_0 <= 16'sh0;
    end else if (_T_46) begin
      adjShiftRegOut_0 <= io_in_bits;
    end
    if (reset) begin
      adjShiftRegOut_1 <= 16'sh0;
    end else if (_T_45) begin
      adjShiftRegOut_1 <= adjShiftRegOut_0;
    end
    if (reset) begin
      adjShiftRegOut_2 <= 16'sh0;
    end else if (_T_44) begin
      adjShiftRegOut_2 <= adjShiftRegOut_1;
    end
    if (reset) begin
      adjShiftRegOut_3 <= 16'sh0;
    end else if (_T_43) begin
      adjShiftRegOut_3 <= adjShiftRegOut_2;
    end
    if (reset) begin
      adjShiftRegOut_4 <= 16'sh0;
    end else if (_T_42) begin
      adjShiftRegOut_4 <= adjShiftRegOut_3;
    end
    if (reset) begin
      adjShiftRegOut_5 <= 16'sh0;
    end else if (_T_41) begin
      adjShiftRegOut_5 <= adjShiftRegOut_4;
    end
    if (reset) begin
      adjShiftRegOut_6 <= 16'sh0;
    end else if (_T_40) begin
      adjShiftRegOut_6 <= adjShiftRegOut_5;
    end
    if (reset) begin
      adjShiftRegOut_7 <= 16'sh0;
    end else if (_T_39) begin
      adjShiftRegOut_7 <= adjShiftRegOut_6;
    end
    if (reset) begin
      cntIn <= 4'h0;
    end else if (_T_132) begin
      cntIn <= 4'h0;
    end else if (_T_1) begin
      cntIn <= _T_62;
    end
    if (reset) begin
      _T_120 <= 1'h0;
    end else if (_T_73) begin
      _T_120 <= _T_59;
    end
    if (reset) begin
      _T_121 <= 1'h0;
    end else if (_T_118) begin
      _T_121 <= _T_120;
    end
    if (reset) begin
      _T_122 <= 1'h0;
    end else if (_T_117) begin
      _T_122 <= _T_121;
    end
    if (reset) begin
      _T_123 <= 1'h0;
    end else if (_T_116) begin
      _T_123 <= _T_122;
    end
    if (reset) begin
      _T_124 <= 1'h0;
    end else if (_T_115) begin
      _T_124 <= _T_123;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else if (_T_114) begin
      _T_125 <= _T_124;
    end
    if (reset) begin
      _T_126 <= 1'h0;
    end else if (_T_113) begin
      _T_126 <= _T_125;
    end
    if (reset) begin
      _T_127 <= 1'h0;
    end else if (_T_112) begin
      _T_127 <= _T_126;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:345 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 345:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[CFARUtils.scala 345:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:330 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 330:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[CFARUtils.scala 330:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CellUnderTest(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut
);
  reg  initialInDone; // @[CFARUtils.scala 453:30]
  reg [31:0] _RAND_0;
  reg  last; // @[CFARUtils.scala 455:21]
  reg [31:0] _RAND_1;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[CFARUtils.scala 457:25]
  wire  _T_3; // @[CFARUtils.scala 457:22]
  wire  _GEN_0; // @[CFARUtils.scala 457:41]
  wire  _T_5; // @[CFARUtils.scala 461:34]
  wire  en; // @[CFARUtils.scala 461:25]
  reg [15:0] cut; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  wire  _T_7; // @[CFARUtils.scala 468:19]
  wire  _GEN_2; // @[CFARUtils.scala 468:36]
  reg  lastOut; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  wire  _T_9; // @[CFARUtils.scala 475:17]
  wire  _T_11; // @[CFARUtils.scala 480:55]
  wire  _T_12; // @[CFARUtils.scala 480:52]
  wire  _T_14; // @[CFARUtils.scala 483:35]
  wire  _T_15; // @[CFARUtils.scala 483:59]
  assign _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = ~initialInDone; // @[CFARUtils.scala 457:25]
  assign _T_3 = _T_1 & _T_2; // @[CFARUtils.scala 457:22]
  assign _GEN_0 = _T_3 | initialInDone; // @[CFARUtils.scala 457:41]
  assign _T_5 = last & io_out_ready; // @[CFARUtils.scala 461:34]
  assign en = _T_1 | _T_5; // @[CFARUtils.scala 461:25]
  assign _T_7 = io_lastIn & _T_1; // @[CFARUtils.scala 468:19]
  assign _GEN_2 = _T_7 | last; // @[CFARUtils.scala 468:36]
  assign _T_9 = lastOut & io_out_ready; // @[CFARUtils.scala 475:17]
  assign _T_11 = ~last; // @[CFARUtils.scala 480:55]
  assign _T_12 = io_out_ready & _T_11; // @[CFARUtils.scala 480:52]
  assign _T_14 = initialInDone & io_in_valid; // @[CFARUtils.scala 483:35]
  assign _T_15 = last & en; // @[CFARUtils.scala 483:59]
  assign io_in_ready = _T_2 | _T_12; // @[CFARUtils.scala 480:18]
  assign io_out_valid = _T_14 | _T_15; // @[CFARUtils.scala 483:18]
  assign io_out_bits = cut; // @[CFARUtils.scala 481:18]
  assign io_lastOut = lastOut; // @[CFARUtils.scala 482:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  initialInDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  last = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cut = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  lastOut = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      initialInDone <= 1'h0;
    end else if (_T_9) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_0;
    end
    if (reset) begin
      last <= 1'h0;
    end else if (_T_9) begin
      last <= 1'h0;
    end else begin
      last <= _GEN_2;
    end
    if (reset) begin
      cut <= 16'sh0;
    end else if (en) begin
      cut <= io_in_bits;
    end
    if (reset) begin
      lastOut <= 1'h0;
    end else if (io_out_ready) begin
      lastOut <= _T_7;
    end
  end
endmodule
module AdjustableShiftRegisterStream_3(
  input         clock,
  input         reset,
  input  [6:0]  io_depth,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_parallelOut_0,
  output [15:0] io_parallelOut_1,
  output [15:0] io_parallelOut_2,
  output [15:0] io_parallelOut_3,
  output [15:0] io_parallelOut_4,
  output [15:0] io_parallelOut_5,
  output [15:0] io_parallelOut_6,
  output [15:0] io_parallelOut_7,
  output [15:0] io_parallelOut_8,
  output [15:0] io_parallelOut_9,
  output [15:0] io_parallelOut_10,
  output [15:0] io_parallelOut_11,
  output [15:0] io_parallelOut_12,
  output [15:0] io_parallelOut_13,
  output [15:0] io_parallelOut_14,
  output [15:0] io_parallelOut_15,
  output [15:0] io_parallelOut_16,
  output [15:0] io_parallelOut_17,
  output [15:0] io_parallelOut_18,
  output [15:0] io_parallelOut_19,
  output [15:0] io_parallelOut_20,
  output [15:0] io_parallelOut_21,
  output [15:0] io_parallelOut_22,
  output [15:0] io_parallelOut_23,
  output [15:0] io_parallelOut_24,
  output [15:0] io_parallelOut_25,
  output [15:0] io_parallelOut_26,
  output [15:0] io_parallelOut_27,
  output [15:0] io_parallelOut_28,
  output [15:0] io_parallelOut_29,
  output [15:0] io_parallelOut_30,
  output [15:0] io_parallelOut_31,
  output [15:0] io_parallelOut_32,
  output [15:0] io_parallelOut_33,
  output [15:0] io_parallelOut_34,
  output [15:0] io_parallelOut_35,
  output [15:0] io_parallelOut_36,
  output [15:0] io_parallelOut_37,
  output [15:0] io_parallelOut_38,
  output [15:0] io_parallelOut_39,
  output [15:0] io_parallelOut_40,
  output [15:0] io_parallelOut_41,
  output [15:0] io_parallelOut_42,
  output [15:0] io_parallelOut_43,
  output [15:0] io_parallelOut_44,
  output [15:0] io_parallelOut_45,
  output [15:0] io_parallelOut_46,
  output [15:0] io_parallelOut_47,
  output [15:0] io_parallelOut_48,
  output [15:0] io_parallelOut_49,
  output [15:0] io_parallelOut_50,
  output [15:0] io_parallelOut_51,
  output [15:0] io_parallelOut_52,
  output [15:0] io_parallelOut_53,
  output [15:0] io_parallelOut_54,
  output [15:0] io_parallelOut_55,
  output [15:0] io_parallelOut_56,
  output [15:0] io_parallelOut_57,
  output [15:0] io_parallelOut_58,
  output [15:0] io_parallelOut_59,
  output [15:0] io_parallelOut_60,
  output [15:0] io_parallelOut_61,
  output [15:0] io_parallelOut_62,
  output [15:0] io_parallelOut_63,
  output [6:0]  io_cnt,
  output        io_regFull
);
  reg  InitialInDone; // @[CFARUtils.scala 379:30]
  reg [31:0] _RAND_0;
  reg  last; // @[CFARUtils.scala 380:21]
  reg [31:0] _RAND_1;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[CFARUtils.scala 385:34]
  wire  en; // @[CFARUtils.scala 385:25]
  wire  _T_3; // @[CFARUtils.scala 345:18]
  wire  _T_5; // @[CFARUtils.scala 345:11]
  wire  _T_6; // @[CFARUtils.scala 345:11]
  wire [6:0] _T_8; // @[CFARUtils.scala 350:87]
  wire  _T_9; // @[CFARUtils.scala 350:78]
  wire  _T_13; // @[CFARUtils.scala 350:78]
  wire  _T_14; // @[CFARUtils.scala 350:94]
  wire  _T_17; // @[CFARUtils.scala 350:78]
  wire  _T_18; // @[CFARUtils.scala 350:94]
  wire  _T_21; // @[CFARUtils.scala 350:78]
  wire  _T_22; // @[CFARUtils.scala 350:94]
  wire  _T_25; // @[CFARUtils.scala 350:78]
  wire  _T_26; // @[CFARUtils.scala 350:94]
  wire  _T_29; // @[CFARUtils.scala 350:78]
  wire  _T_30; // @[CFARUtils.scala 350:94]
  wire  _T_33; // @[CFARUtils.scala 350:78]
  wire  _T_34; // @[CFARUtils.scala 350:94]
  wire  _T_37; // @[CFARUtils.scala 350:78]
  wire  _T_38; // @[CFARUtils.scala 350:94]
  wire  _T_41; // @[CFARUtils.scala 350:78]
  wire  _T_42; // @[CFARUtils.scala 350:94]
  wire  _T_45; // @[CFARUtils.scala 350:78]
  wire  _T_46; // @[CFARUtils.scala 350:94]
  wire  _T_49; // @[CFARUtils.scala 350:78]
  wire  _T_50; // @[CFARUtils.scala 350:94]
  wire  _T_53; // @[CFARUtils.scala 350:78]
  wire  _T_54; // @[CFARUtils.scala 350:94]
  wire  _T_57; // @[CFARUtils.scala 350:78]
  wire  _T_58; // @[CFARUtils.scala 350:94]
  wire  _T_61; // @[CFARUtils.scala 350:78]
  wire  _T_62; // @[CFARUtils.scala 350:94]
  wire  _T_65; // @[CFARUtils.scala 350:78]
  wire  _T_66; // @[CFARUtils.scala 350:94]
  wire  _T_69; // @[CFARUtils.scala 350:78]
  wire  _T_70; // @[CFARUtils.scala 350:94]
  wire  _T_73; // @[CFARUtils.scala 350:78]
  wire  _T_74; // @[CFARUtils.scala 350:94]
  wire  _T_77; // @[CFARUtils.scala 350:78]
  wire  _T_78; // @[CFARUtils.scala 350:94]
  wire  _T_81; // @[CFARUtils.scala 350:78]
  wire  _T_82; // @[CFARUtils.scala 350:94]
  wire  _T_85; // @[CFARUtils.scala 350:78]
  wire  _T_86; // @[CFARUtils.scala 350:94]
  wire  _T_89; // @[CFARUtils.scala 350:78]
  wire  _T_90; // @[CFARUtils.scala 350:94]
  wire  _T_93; // @[CFARUtils.scala 350:78]
  wire  _T_94; // @[CFARUtils.scala 350:94]
  wire  _T_97; // @[CFARUtils.scala 350:78]
  wire  _T_98; // @[CFARUtils.scala 350:94]
  wire  _T_101; // @[CFARUtils.scala 350:78]
  wire  _T_102; // @[CFARUtils.scala 350:94]
  wire  _T_105; // @[CFARUtils.scala 350:78]
  wire  _T_106; // @[CFARUtils.scala 350:94]
  wire  _T_109; // @[CFARUtils.scala 350:78]
  wire  _T_110; // @[CFARUtils.scala 350:94]
  wire  _T_113; // @[CFARUtils.scala 350:78]
  wire  _T_114; // @[CFARUtils.scala 350:94]
  wire  _T_117; // @[CFARUtils.scala 350:78]
  wire  _T_118; // @[CFARUtils.scala 350:94]
  wire  _T_121; // @[CFARUtils.scala 350:78]
  wire  _T_122; // @[CFARUtils.scala 350:94]
  wire  _T_125; // @[CFARUtils.scala 350:78]
  wire  _T_126; // @[CFARUtils.scala 350:94]
  wire  _T_129; // @[CFARUtils.scala 350:78]
  wire  _T_130; // @[CFARUtils.scala 350:94]
  wire  _T_133; // @[CFARUtils.scala 350:78]
  wire  _T_134; // @[CFARUtils.scala 350:94]
  wire  _T_137; // @[CFARUtils.scala 350:78]
  wire  _T_138; // @[CFARUtils.scala 350:94]
  wire  _T_141; // @[CFARUtils.scala 350:78]
  wire  _T_142; // @[CFARUtils.scala 350:94]
  wire  _T_145; // @[CFARUtils.scala 350:78]
  wire  _T_146; // @[CFARUtils.scala 350:94]
  wire  _T_149; // @[CFARUtils.scala 350:78]
  wire  _T_150; // @[CFARUtils.scala 350:94]
  wire  _T_153; // @[CFARUtils.scala 350:78]
  wire  _T_154; // @[CFARUtils.scala 350:94]
  wire  _T_157; // @[CFARUtils.scala 350:78]
  wire  _T_158; // @[CFARUtils.scala 350:94]
  wire  _T_161; // @[CFARUtils.scala 350:78]
  wire  _T_162; // @[CFARUtils.scala 350:94]
  wire  _T_165; // @[CFARUtils.scala 350:78]
  wire  _T_166; // @[CFARUtils.scala 350:94]
  wire  _T_169; // @[CFARUtils.scala 350:78]
  wire  _T_170; // @[CFARUtils.scala 350:94]
  wire  _T_173; // @[CFARUtils.scala 350:78]
  wire  _T_174; // @[CFARUtils.scala 350:94]
  wire  _T_177; // @[CFARUtils.scala 350:78]
  wire  _T_178; // @[CFARUtils.scala 350:94]
  wire  _T_181; // @[CFARUtils.scala 350:78]
  wire  _T_182; // @[CFARUtils.scala 350:94]
  wire  _T_185; // @[CFARUtils.scala 350:78]
  wire  _T_186; // @[CFARUtils.scala 350:94]
  wire  _T_189; // @[CFARUtils.scala 350:78]
  wire  _T_190; // @[CFARUtils.scala 350:94]
  wire  _T_193; // @[CFARUtils.scala 350:78]
  wire  _T_194; // @[CFARUtils.scala 350:94]
  wire  _T_197; // @[CFARUtils.scala 350:78]
  wire  _T_198; // @[CFARUtils.scala 350:94]
  wire  _T_201; // @[CFARUtils.scala 350:78]
  wire  _T_202; // @[CFARUtils.scala 350:94]
  wire  _T_205; // @[CFARUtils.scala 350:78]
  wire  _T_206; // @[CFARUtils.scala 350:94]
  wire  _T_209; // @[CFARUtils.scala 350:78]
  wire  _T_210; // @[CFARUtils.scala 350:94]
  wire  _T_213; // @[CFARUtils.scala 350:78]
  wire  _T_214; // @[CFARUtils.scala 350:94]
  wire  _T_217; // @[CFARUtils.scala 350:78]
  wire  _T_218; // @[CFARUtils.scala 350:94]
  wire  _T_221; // @[CFARUtils.scala 350:78]
  wire  _T_222; // @[CFARUtils.scala 350:94]
  wire  _T_225; // @[CFARUtils.scala 350:78]
  wire  _T_226; // @[CFARUtils.scala 350:94]
  wire  _T_229; // @[CFARUtils.scala 350:78]
  wire  _T_230; // @[CFARUtils.scala 350:94]
  wire  _T_233; // @[CFARUtils.scala 350:78]
  wire  _T_234; // @[CFARUtils.scala 350:94]
  wire  _T_237; // @[CFARUtils.scala 350:78]
  wire  _T_238; // @[CFARUtils.scala 350:94]
  wire  _T_241; // @[CFARUtils.scala 350:78]
  wire  _T_242; // @[CFARUtils.scala 350:94]
  wire  _T_245; // @[CFARUtils.scala 350:78]
  wire  _T_246; // @[CFARUtils.scala 350:94]
  wire  _T_249; // @[CFARUtils.scala 350:78]
  wire  _T_250; // @[CFARUtils.scala 350:94]
  wire  _T_253; // @[CFARUtils.scala 350:78]
  wire  _T_254; // @[CFARUtils.scala 350:94]
  wire  _T_257; // @[CFARUtils.scala 350:78]
  wire  _T_258; // @[CFARUtils.scala 350:94]
  wire  _T_261; // @[CFARUtils.scala 350:78]
  wire  _T_262; // @[CFARUtils.scala 350:94]
  wire  activeRegs_63; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_263; // @[CFARUtils.scala 319:37]
  wire  activeRegs_62; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_264; // @[CFARUtils.scala 319:37]
  wire  activeRegs_61; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_265; // @[CFARUtils.scala 319:37]
  wire  activeRegs_60; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_266; // @[CFARUtils.scala 319:37]
  wire  activeRegs_59; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_267; // @[CFARUtils.scala 319:37]
  wire  activeRegs_58; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_268; // @[CFARUtils.scala 319:37]
  wire  activeRegs_57; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_269; // @[CFARUtils.scala 319:37]
  wire  activeRegs_56; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_270; // @[CFARUtils.scala 319:37]
  wire  activeRegs_55; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_271; // @[CFARUtils.scala 319:37]
  wire  activeRegs_54; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_272; // @[CFARUtils.scala 319:37]
  wire  activeRegs_53; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_273; // @[CFARUtils.scala 319:37]
  wire  activeRegs_52; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_274; // @[CFARUtils.scala 319:37]
  wire  activeRegs_51; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_275; // @[CFARUtils.scala 319:37]
  wire  activeRegs_50; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_276; // @[CFARUtils.scala 319:37]
  wire  activeRegs_49; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_277; // @[CFARUtils.scala 319:37]
  wire  activeRegs_48; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_278; // @[CFARUtils.scala 319:37]
  wire  activeRegs_47; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_279; // @[CFARUtils.scala 319:37]
  wire  activeRegs_46; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_280; // @[CFARUtils.scala 319:37]
  wire  activeRegs_45; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_281; // @[CFARUtils.scala 319:37]
  wire  activeRegs_44; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_282; // @[CFARUtils.scala 319:37]
  wire  activeRegs_43; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_283; // @[CFARUtils.scala 319:37]
  wire  activeRegs_42; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_284; // @[CFARUtils.scala 319:37]
  wire  activeRegs_41; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_285; // @[CFARUtils.scala 319:37]
  wire  activeRegs_40; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_286; // @[CFARUtils.scala 319:37]
  wire  activeRegs_39; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_287; // @[CFARUtils.scala 319:37]
  wire  activeRegs_38; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_288; // @[CFARUtils.scala 319:37]
  wire  activeRegs_37; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_289; // @[CFARUtils.scala 319:37]
  wire  activeRegs_36; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_290; // @[CFARUtils.scala 319:37]
  wire  activeRegs_35; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_291; // @[CFARUtils.scala 319:37]
  wire  activeRegs_34; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_292; // @[CFARUtils.scala 319:37]
  wire  activeRegs_33; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_293; // @[CFARUtils.scala 319:37]
  wire  activeRegs_32; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_294; // @[CFARUtils.scala 319:37]
  wire  activeRegs_31; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_295; // @[CFARUtils.scala 319:37]
  wire  activeRegs_30; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_296; // @[CFARUtils.scala 319:37]
  wire  activeRegs_29; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_297; // @[CFARUtils.scala 319:37]
  wire  activeRegs_28; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_298; // @[CFARUtils.scala 319:37]
  wire  activeRegs_27; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_299; // @[CFARUtils.scala 319:37]
  wire  activeRegs_26; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_300; // @[CFARUtils.scala 319:37]
  wire  activeRegs_25; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_301; // @[CFARUtils.scala 319:37]
  wire  activeRegs_24; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_302; // @[CFARUtils.scala 319:37]
  wire  activeRegs_23; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_303; // @[CFARUtils.scala 319:37]
  wire  activeRegs_22; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_304; // @[CFARUtils.scala 319:37]
  wire  activeRegs_21; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_305; // @[CFARUtils.scala 319:37]
  wire  activeRegs_20; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_306; // @[CFARUtils.scala 319:37]
  wire  activeRegs_19; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_307; // @[CFARUtils.scala 319:37]
  wire  activeRegs_18; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_308; // @[CFARUtils.scala 319:37]
  wire  activeRegs_17; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_309; // @[CFARUtils.scala 319:37]
  wire  activeRegs_16; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_310; // @[CFARUtils.scala 319:37]
  wire  activeRegs_15; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_311; // @[CFARUtils.scala 319:37]
  wire  activeRegs_14; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_312; // @[CFARUtils.scala 319:37]
  wire  activeRegs_13; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_313; // @[CFARUtils.scala 319:37]
  wire  activeRegs_12; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_314; // @[CFARUtils.scala 319:37]
  wire  activeRegs_11; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_315; // @[CFARUtils.scala 319:37]
  wire  activeRegs_10; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_316; // @[CFARUtils.scala 319:37]
  wire  activeRegs_9; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_317; // @[CFARUtils.scala 319:37]
  wire  activeRegs_8; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_318; // @[CFARUtils.scala 319:37]
  wire  activeRegs_7; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_319; // @[CFARUtils.scala 319:37]
  wire  activeRegs_6; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_320; // @[CFARUtils.scala 319:37]
  wire  activeRegs_5; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_321; // @[CFARUtils.scala 319:37]
  wire  activeRegs_4; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_322; // @[CFARUtils.scala 319:37]
  wire  activeRegs_3; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_323; // @[CFARUtils.scala 319:37]
  wire  activeRegs_2; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_324; // @[CFARUtils.scala 319:37]
  wire  activeRegs_1; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_325; // @[CFARUtils.scala 319:37]
  wire  activeRegs_0; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  wire  _T_326; // @[CFARUtils.scala 319:37]
  reg [15:0] adjShiftRegOut_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [15:0] adjShiftRegOut_1; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [15:0] adjShiftRegOut_2; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [15:0] adjShiftRegOut_3; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [15:0] adjShiftRegOut_4; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [15:0] adjShiftRegOut_5; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [15:0] adjShiftRegOut_6; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  reg [15:0] adjShiftRegOut_7; // @[Reg.scala 27:20]
  reg [31:0] _RAND_9;
  reg [15:0] adjShiftRegOut_8; // @[Reg.scala 27:20]
  reg [31:0] _RAND_10;
  reg [15:0] adjShiftRegOut_9; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg [15:0] adjShiftRegOut_10; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg [15:0] adjShiftRegOut_11; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg [15:0] adjShiftRegOut_12; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  reg [15:0] adjShiftRegOut_13; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  reg [15:0] adjShiftRegOut_14; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg [15:0] adjShiftRegOut_15; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  reg [15:0] adjShiftRegOut_16; // @[Reg.scala 27:20]
  reg [31:0] _RAND_18;
  reg [15:0] adjShiftRegOut_17; // @[Reg.scala 27:20]
  reg [31:0] _RAND_19;
  reg [15:0] adjShiftRegOut_18; // @[Reg.scala 27:20]
  reg [31:0] _RAND_20;
  reg [15:0] adjShiftRegOut_19; // @[Reg.scala 27:20]
  reg [31:0] _RAND_21;
  reg [15:0] adjShiftRegOut_20; // @[Reg.scala 27:20]
  reg [31:0] _RAND_22;
  reg [15:0] adjShiftRegOut_21; // @[Reg.scala 27:20]
  reg [31:0] _RAND_23;
  reg [15:0] adjShiftRegOut_22; // @[Reg.scala 27:20]
  reg [31:0] _RAND_24;
  reg [15:0] adjShiftRegOut_23; // @[Reg.scala 27:20]
  reg [31:0] _RAND_25;
  reg [15:0] adjShiftRegOut_24; // @[Reg.scala 27:20]
  reg [31:0] _RAND_26;
  reg [15:0] adjShiftRegOut_25; // @[Reg.scala 27:20]
  reg [31:0] _RAND_27;
  reg [15:0] adjShiftRegOut_26; // @[Reg.scala 27:20]
  reg [31:0] _RAND_28;
  reg [15:0] adjShiftRegOut_27; // @[Reg.scala 27:20]
  reg [31:0] _RAND_29;
  reg [15:0] adjShiftRegOut_28; // @[Reg.scala 27:20]
  reg [31:0] _RAND_30;
  reg [15:0] adjShiftRegOut_29; // @[Reg.scala 27:20]
  reg [31:0] _RAND_31;
  reg [15:0] adjShiftRegOut_30; // @[Reg.scala 27:20]
  reg [31:0] _RAND_32;
  reg [15:0] adjShiftRegOut_31; // @[Reg.scala 27:20]
  reg [31:0] _RAND_33;
  reg [15:0] adjShiftRegOut_32; // @[Reg.scala 27:20]
  reg [31:0] _RAND_34;
  reg [15:0] adjShiftRegOut_33; // @[Reg.scala 27:20]
  reg [31:0] _RAND_35;
  reg [15:0] adjShiftRegOut_34; // @[Reg.scala 27:20]
  reg [31:0] _RAND_36;
  reg [15:0] adjShiftRegOut_35; // @[Reg.scala 27:20]
  reg [31:0] _RAND_37;
  reg [15:0] adjShiftRegOut_36; // @[Reg.scala 27:20]
  reg [31:0] _RAND_38;
  reg [15:0] adjShiftRegOut_37; // @[Reg.scala 27:20]
  reg [31:0] _RAND_39;
  reg [15:0] adjShiftRegOut_38; // @[Reg.scala 27:20]
  reg [31:0] _RAND_40;
  reg [15:0] adjShiftRegOut_39; // @[Reg.scala 27:20]
  reg [31:0] _RAND_41;
  reg [15:0] adjShiftRegOut_40; // @[Reg.scala 27:20]
  reg [31:0] _RAND_42;
  reg [15:0] adjShiftRegOut_41; // @[Reg.scala 27:20]
  reg [31:0] _RAND_43;
  reg [15:0] adjShiftRegOut_42; // @[Reg.scala 27:20]
  reg [31:0] _RAND_44;
  reg [15:0] adjShiftRegOut_43; // @[Reg.scala 27:20]
  reg [31:0] _RAND_45;
  reg [15:0] adjShiftRegOut_44; // @[Reg.scala 27:20]
  reg [31:0] _RAND_46;
  reg [15:0] adjShiftRegOut_45; // @[Reg.scala 27:20]
  reg [31:0] _RAND_47;
  reg [15:0] adjShiftRegOut_46; // @[Reg.scala 27:20]
  reg [31:0] _RAND_48;
  reg [15:0] adjShiftRegOut_47; // @[Reg.scala 27:20]
  reg [31:0] _RAND_49;
  reg [15:0] adjShiftRegOut_48; // @[Reg.scala 27:20]
  reg [31:0] _RAND_50;
  reg [15:0] adjShiftRegOut_49; // @[Reg.scala 27:20]
  reg [31:0] _RAND_51;
  reg [15:0] adjShiftRegOut_50; // @[Reg.scala 27:20]
  reg [31:0] _RAND_52;
  reg [15:0] adjShiftRegOut_51; // @[Reg.scala 27:20]
  reg [31:0] _RAND_53;
  reg [15:0] adjShiftRegOut_52; // @[Reg.scala 27:20]
  reg [31:0] _RAND_54;
  reg [15:0] adjShiftRegOut_53; // @[Reg.scala 27:20]
  reg [31:0] _RAND_55;
  reg [15:0] adjShiftRegOut_54; // @[Reg.scala 27:20]
  reg [31:0] _RAND_56;
  reg [15:0] adjShiftRegOut_55; // @[Reg.scala 27:20]
  reg [31:0] _RAND_57;
  reg [15:0] adjShiftRegOut_56; // @[Reg.scala 27:20]
  reg [31:0] _RAND_58;
  reg [15:0] adjShiftRegOut_57; // @[Reg.scala 27:20]
  reg [31:0] _RAND_59;
  reg [15:0] adjShiftRegOut_58; // @[Reg.scala 27:20]
  reg [31:0] _RAND_60;
  reg [15:0] adjShiftRegOut_59; // @[Reg.scala 27:20]
  reg [31:0] _RAND_61;
  reg [15:0] adjShiftRegOut_60; // @[Reg.scala 27:20]
  reg [31:0] _RAND_62;
  reg [15:0] adjShiftRegOut_61; // @[Reg.scala 27:20]
  reg [31:0] _RAND_63;
  reg [15:0] adjShiftRegOut_62; // @[Reg.scala 27:20]
  reg [31:0] _RAND_64;
  reg [15:0] adjShiftRegOut_63; // @[Reg.scala 27:20]
  reg [31:0] _RAND_65;
  reg [6:0] cntIn; // @[CFARUtils.scala 390:23]
  reg [31:0] _RAND_66;
  wire  _T_395; // @[CFARUtils.scala 392:19]
  wire  _GEN_64; // @[CFARUtils.scala 392:36]
  wire [6:0] _T_398; // @[CFARUtils.scala 397:20]
  wire  _T_399; // @[CFARUtils.scala 400:18]
  wire  _T_402; // @[CFARUtils.scala 401:17]
  wire  _T_404; // @[CFARUtils.scala 401:36]
  wire  _GEN_66; // @[CFARUtils.scala 401:53]
  wire  _T_406; // @[CFARUtils.scala 406:36]
  wire  _T_407; // @[CFARUtils.scala 406:24]
  wire  _GEN_67; // @[CFARUtils.scala 406:45]
  wire  _T_409; // @[Decoupled.scala 40:37]
  wire  _T_672; // @[CFARUtils.scala 319:37]
  wire  _T_673; // @[CFARUtils.scala 319:37]
  wire  _T_674; // @[CFARUtils.scala 319:37]
  wire  _T_675; // @[CFARUtils.scala 319:37]
  wire  _T_676; // @[CFARUtils.scala 319:37]
  wire  _T_677; // @[CFARUtils.scala 319:37]
  wire  _T_678; // @[CFARUtils.scala 319:37]
  wire  _T_679; // @[CFARUtils.scala 319:37]
  wire  _T_680; // @[CFARUtils.scala 319:37]
  wire  _T_681; // @[CFARUtils.scala 319:37]
  wire  _T_682; // @[CFARUtils.scala 319:37]
  wire  _T_683; // @[CFARUtils.scala 319:37]
  wire  _T_684; // @[CFARUtils.scala 319:37]
  wire  _T_685; // @[CFARUtils.scala 319:37]
  wire  _T_686; // @[CFARUtils.scala 319:37]
  wire  _T_687; // @[CFARUtils.scala 319:37]
  wire  _T_688; // @[CFARUtils.scala 319:37]
  wire  _T_689; // @[CFARUtils.scala 319:37]
  wire  _T_690; // @[CFARUtils.scala 319:37]
  wire  _T_691; // @[CFARUtils.scala 319:37]
  wire  _T_692; // @[CFARUtils.scala 319:37]
  wire  _T_693; // @[CFARUtils.scala 319:37]
  wire  _T_694; // @[CFARUtils.scala 319:37]
  wire  _T_695; // @[CFARUtils.scala 319:37]
  wire  _T_696; // @[CFARUtils.scala 319:37]
  wire  _T_697; // @[CFARUtils.scala 319:37]
  wire  _T_698; // @[CFARUtils.scala 319:37]
  wire  _T_699; // @[CFARUtils.scala 319:37]
  wire  _T_700; // @[CFARUtils.scala 319:37]
  wire  _T_701; // @[CFARUtils.scala 319:37]
  wire  _T_702; // @[CFARUtils.scala 319:37]
  wire  _T_703; // @[CFARUtils.scala 319:37]
  wire  _T_704; // @[CFARUtils.scala 319:37]
  wire  _T_705; // @[CFARUtils.scala 319:37]
  wire  _T_706; // @[CFARUtils.scala 319:37]
  wire  _T_707; // @[CFARUtils.scala 319:37]
  wire  _T_708; // @[CFARUtils.scala 319:37]
  wire  _T_709; // @[CFARUtils.scala 319:37]
  wire  _T_710; // @[CFARUtils.scala 319:37]
  wire  _T_711; // @[CFARUtils.scala 319:37]
  wire  _T_712; // @[CFARUtils.scala 319:37]
  wire  _T_713; // @[CFARUtils.scala 319:37]
  wire  _T_714; // @[CFARUtils.scala 319:37]
  wire  _T_715; // @[CFARUtils.scala 319:37]
  wire  _T_716; // @[CFARUtils.scala 319:37]
  wire  _T_717; // @[CFARUtils.scala 319:37]
  wire  _T_718; // @[CFARUtils.scala 319:37]
  wire  _T_719; // @[CFARUtils.scala 319:37]
  wire  _T_720; // @[CFARUtils.scala 319:37]
  wire  _T_721; // @[CFARUtils.scala 319:37]
  wire  _T_722; // @[CFARUtils.scala 319:37]
  wire  _T_723; // @[CFARUtils.scala 319:37]
  wire  _T_724; // @[CFARUtils.scala 319:37]
  wire  _T_725; // @[CFARUtils.scala 319:37]
  wire  _T_726; // @[CFARUtils.scala 319:37]
  wire  _T_727; // @[CFARUtils.scala 319:37]
  wire  _T_728; // @[CFARUtils.scala 319:37]
  wire  _T_729; // @[CFARUtils.scala 319:37]
  wire  _T_730; // @[CFARUtils.scala 319:37]
  wire  _T_731; // @[CFARUtils.scala 319:37]
  wire  _T_732; // @[CFARUtils.scala 319:37]
  wire  _T_733; // @[CFARUtils.scala 319:37]
  wire  _T_734; // @[CFARUtils.scala 319:37]
  reg  _T_736; // @[Reg.scala 27:20]
  reg [31:0] _RAND_67;
  reg  _T_737; // @[Reg.scala 27:20]
  reg [31:0] _RAND_68;
  reg  _T_738; // @[Reg.scala 27:20]
  reg [31:0] _RAND_69;
  reg  _T_739; // @[Reg.scala 27:20]
  reg [31:0] _RAND_70;
  reg  _T_740; // @[Reg.scala 27:20]
  reg [31:0] _RAND_71;
  reg  _T_741; // @[Reg.scala 27:20]
  reg [31:0] _RAND_72;
  reg  _T_742; // @[Reg.scala 27:20]
  reg [31:0] _RAND_73;
  reg  _T_743; // @[Reg.scala 27:20]
  reg [31:0] _RAND_74;
  reg  _T_744; // @[Reg.scala 27:20]
  reg [31:0] _RAND_75;
  reg  _T_745; // @[Reg.scala 27:20]
  reg [31:0] _RAND_76;
  reg  _T_746; // @[Reg.scala 27:20]
  reg [31:0] _RAND_77;
  reg  _T_747; // @[Reg.scala 27:20]
  reg [31:0] _RAND_78;
  reg  _T_748; // @[Reg.scala 27:20]
  reg [31:0] _RAND_79;
  reg  _T_749; // @[Reg.scala 27:20]
  reg [31:0] _RAND_80;
  reg  _T_750; // @[Reg.scala 27:20]
  reg [31:0] _RAND_81;
  reg  _T_751; // @[Reg.scala 27:20]
  reg [31:0] _RAND_82;
  reg  _T_752; // @[Reg.scala 27:20]
  reg [31:0] _RAND_83;
  reg  _T_753; // @[Reg.scala 27:20]
  reg [31:0] _RAND_84;
  reg  _T_754; // @[Reg.scala 27:20]
  reg [31:0] _RAND_85;
  reg  _T_755; // @[Reg.scala 27:20]
  reg [31:0] _RAND_86;
  reg  _T_756; // @[Reg.scala 27:20]
  reg [31:0] _RAND_87;
  reg  _T_757; // @[Reg.scala 27:20]
  reg [31:0] _RAND_88;
  reg  _T_758; // @[Reg.scala 27:20]
  reg [31:0] _RAND_89;
  reg  _T_759; // @[Reg.scala 27:20]
  reg [31:0] _RAND_90;
  reg  _T_760; // @[Reg.scala 27:20]
  reg [31:0] _RAND_91;
  reg  _T_761; // @[Reg.scala 27:20]
  reg [31:0] _RAND_92;
  reg  _T_762; // @[Reg.scala 27:20]
  reg [31:0] _RAND_93;
  reg  _T_763; // @[Reg.scala 27:20]
  reg [31:0] _RAND_94;
  reg  _T_764; // @[Reg.scala 27:20]
  reg [31:0] _RAND_95;
  reg  _T_765; // @[Reg.scala 27:20]
  reg [31:0] _RAND_96;
  reg  _T_766; // @[Reg.scala 27:20]
  reg [31:0] _RAND_97;
  reg  _T_767; // @[Reg.scala 27:20]
  reg [31:0] _RAND_98;
  reg  _T_768; // @[Reg.scala 27:20]
  reg [31:0] _RAND_99;
  reg  _T_769; // @[Reg.scala 27:20]
  reg [31:0] _RAND_100;
  reg  _T_770; // @[Reg.scala 27:20]
  reg [31:0] _RAND_101;
  reg  _T_771; // @[Reg.scala 27:20]
  reg [31:0] _RAND_102;
  reg  _T_772; // @[Reg.scala 27:20]
  reg [31:0] _RAND_103;
  reg  _T_773; // @[Reg.scala 27:20]
  reg [31:0] _RAND_104;
  reg  _T_774; // @[Reg.scala 27:20]
  reg [31:0] _RAND_105;
  reg  _T_775; // @[Reg.scala 27:20]
  reg [31:0] _RAND_106;
  reg  _T_776; // @[Reg.scala 27:20]
  reg [31:0] _RAND_107;
  reg  _T_777; // @[Reg.scala 27:20]
  reg [31:0] _RAND_108;
  reg  _T_778; // @[Reg.scala 27:20]
  reg [31:0] _RAND_109;
  reg  _T_779; // @[Reg.scala 27:20]
  reg [31:0] _RAND_110;
  reg  _T_780; // @[Reg.scala 27:20]
  reg [31:0] _RAND_111;
  reg  _T_781; // @[Reg.scala 27:20]
  reg [31:0] _RAND_112;
  reg  _T_782; // @[Reg.scala 27:20]
  reg [31:0] _RAND_113;
  reg  _T_783; // @[Reg.scala 27:20]
  reg [31:0] _RAND_114;
  reg  _T_784; // @[Reg.scala 27:20]
  reg [31:0] _RAND_115;
  reg  _T_785; // @[Reg.scala 27:20]
  reg [31:0] _RAND_116;
  reg  _T_786; // @[Reg.scala 27:20]
  reg [31:0] _RAND_117;
  reg  _T_787; // @[Reg.scala 27:20]
  reg [31:0] _RAND_118;
  reg  _T_788; // @[Reg.scala 27:20]
  reg [31:0] _RAND_119;
  reg  _T_789; // @[Reg.scala 27:20]
  reg [31:0] _RAND_120;
  reg  _T_790; // @[Reg.scala 27:20]
  reg [31:0] _RAND_121;
  reg  _T_791; // @[Reg.scala 27:20]
  reg [31:0] _RAND_122;
  reg  _T_792; // @[Reg.scala 27:20]
  reg [31:0] _RAND_123;
  reg  _T_793; // @[Reg.scala 27:20]
  reg [31:0] _RAND_124;
  reg  _T_794; // @[Reg.scala 27:20]
  reg [31:0] _RAND_125;
  reg  _T_795; // @[Reg.scala 27:20]
  reg [31:0] _RAND_126;
  reg  _T_796; // @[Reg.scala 27:20]
  reg [31:0] _RAND_127;
  reg  _T_797; // @[Reg.scala 27:20]
  reg [31:0] _RAND_128;
  reg  _T_798; // @[Reg.scala 27:20]
  reg [31:0] _RAND_129;
  reg  _T_799; // @[Reg.scala 27:20]
  reg [31:0] _RAND_130;
  wire  _GEN_134; // @[CFARUtils.scala 414:17]
  wire  _GEN_135; // @[CFARUtils.scala 414:17]
  wire  _GEN_136; // @[CFARUtils.scala 414:17]
  wire  _GEN_137; // @[CFARUtils.scala 414:17]
  wire  _GEN_138; // @[CFARUtils.scala 414:17]
  wire  _GEN_139; // @[CFARUtils.scala 414:17]
  wire  _GEN_140; // @[CFARUtils.scala 414:17]
  wire  _GEN_141; // @[CFARUtils.scala 414:17]
  wire  _GEN_142; // @[CFARUtils.scala 414:17]
  wire  _GEN_143; // @[CFARUtils.scala 414:17]
  wire  _GEN_144; // @[CFARUtils.scala 414:17]
  wire  _GEN_145; // @[CFARUtils.scala 414:17]
  wire  _GEN_146; // @[CFARUtils.scala 414:17]
  wire  _GEN_147; // @[CFARUtils.scala 414:17]
  wire  _GEN_148; // @[CFARUtils.scala 414:17]
  wire  _GEN_149; // @[CFARUtils.scala 414:17]
  wire  _GEN_150; // @[CFARUtils.scala 414:17]
  wire  _GEN_151; // @[CFARUtils.scala 414:17]
  wire  _GEN_152; // @[CFARUtils.scala 414:17]
  wire  _GEN_153; // @[CFARUtils.scala 414:17]
  wire  _GEN_154; // @[CFARUtils.scala 414:17]
  wire  _GEN_155; // @[CFARUtils.scala 414:17]
  wire  _GEN_156; // @[CFARUtils.scala 414:17]
  wire  _GEN_157; // @[CFARUtils.scala 414:17]
  wire  _GEN_158; // @[CFARUtils.scala 414:17]
  wire  _GEN_159; // @[CFARUtils.scala 414:17]
  wire  _GEN_160; // @[CFARUtils.scala 414:17]
  wire  _GEN_161; // @[CFARUtils.scala 414:17]
  wire  _GEN_162; // @[CFARUtils.scala 414:17]
  wire  _GEN_163; // @[CFARUtils.scala 414:17]
  wire  _GEN_164; // @[CFARUtils.scala 414:17]
  wire  _GEN_165; // @[CFARUtils.scala 414:17]
  wire  _GEN_166; // @[CFARUtils.scala 414:17]
  wire  _GEN_167; // @[CFARUtils.scala 414:17]
  wire  _GEN_168; // @[CFARUtils.scala 414:17]
  wire  _GEN_169; // @[CFARUtils.scala 414:17]
  wire  _GEN_170; // @[CFARUtils.scala 414:17]
  wire  _GEN_171; // @[CFARUtils.scala 414:17]
  wire  _GEN_172; // @[CFARUtils.scala 414:17]
  wire  _GEN_173; // @[CFARUtils.scala 414:17]
  wire  _GEN_174; // @[CFARUtils.scala 414:17]
  wire  _GEN_175; // @[CFARUtils.scala 414:17]
  wire  _GEN_176; // @[CFARUtils.scala 414:17]
  wire  _GEN_177; // @[CFARUtils.scala 414:17]
  wire  _GEN_178; // @[CFARUtils.scala 414:17]
  wire  _GEN_179; // @[CFARUtils.scala 414:17]
  wire  _GEN_180; // @[CFARUtils.scala 414:17]
  wire  _GEN_181; // @[CFARUtils.scala 414:17]
  wire  _GEN_182; // @[CFARUtils.scala 414:17]
  wire  _GEN_183; // @[CFARUtils.scala 414:17]
  wire  _GEN_184; // @[CFARUtils.scala 414:17]
  wire  _GEN_185; // @[CFARUtils.scala 414:17]
  wire  _GEN_186; // @[CFARUtils.scala 414:17]
  wire  _GEN_187; // @[CFARUtils.scala 414:17]
  wire  _GEN_188; // @[CFARUtils.scala 414:17]
  wire  _GEN_189; // @[CFARUtils.scala 414:17]
  wire  _GEN_190; // @[CFARUtils.scala 414:17]
  wire  _GEN_191; // @[CFARUtils.scala 414:17]
  wire  _GEN_192; // @[CFARUtils.scala 414:17]
  wire  _GEN_193; // @[CFARUtils.scala 414:17]
  wire  _GEN_194; // @[CFARUtils.scala 414:17]
  wire  _GEN_195; // @[CFARUtils.scala 414:17]
  wire  _GEN_196; // @[CFARUtils.scala 414:17]
  wire  _T_804; // @[CFARUtils.scala 414:17]
  wire  _T_808; // @[CFARUtils.scala 421:36]
  wire  _T_810; // @[CFARUtils.scala 429:37]
  wire  _T_812; // @[CFARUtils.scala 429:73]
  wire  _T_821; // @[CFARUtils.scala 436:70]
  wire  _T_822; // @[CFARUtils.scala 436:94]
  wire  _T_823; // @[CFARUtils.scala 436:85]
  assign _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = last & io_out_ready; // @[CFARUtils.scala 385:34]
  assign en = _T_1 | _T_2; // @[CFARUtils.scala 385:25]
  assign _T_3 = io_depth <= 7'h40; // @[CFARUtils.scala 345:18]
  assign _T_5 = _T_3 | reset; // @[CFARUtils.scala 345:11]
  assign _T_6 = ~_T_5; // @[CFARUtils.scala 345:11]
  assign _T_8 = io_depth - 7'h1; // @[CFARUtils.scala 350:87]
  assign _T_9 = 1'h1; // @[CFARUtils.scala 350:78]
  assign _T_13 = 7'h1 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_14 = _T_13; // @[CFARUtils.scala 350:94]
  assign _T_17 = 7'h2 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_18 = _T_17; // @[CFARUtils.scala 350:94]
  assign _T_21 = 7'h3 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_22 = _T_21; // @[CFARUtils.scala 350:94]
  assign _T_25 = 7'h4 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_26 = _T_25; // @[CFARUtils.scala 350:94]
  assign _T_29 = 7'h5 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_30 = _T_29; // @[CFARUtils.scala 350:94]
  assign _T_33 = 7'h6 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_34 = _T_33; // @[CFARUtils.scala 350:94]
  assign _T_37 = 7'h7 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_38 = _T_37; // @[CFARUtils.scala 350:94]
  assign _T_41 = 7'h8 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_42 = _T_41; // @[CFARUtils.scala 350:94]
  assign _T_45 = 7'h9 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_46 = _T_45; // @[CFARUtils.scala 350:94]
  assign _T_49 = 7'ha <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_50 = _T_49; // @[CFARUtils.scala 350:94]
  assign _T_53 = 7'hb <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_54 = _T_53; // @[CFARUtils.scala 350:94]
  assign _T_57 = 7'hc <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_58 = _T_57; // @[CFARUtils.scala 350:94]
  assign _T_61 = 7'hd <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_62 = _T_61; // @[CFARUtils.scala 350:94]
  assign _T_65 = 7'he <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_66 = _T_65; // @[CFARUtils.scala 350:94]
  assign _T_69 = 7'hf <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_70 = _T_69; // @[CFARUtils.scala 350:94]
  assign _T_73 = 7'h10 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_74 = _T_73; // @[CFARUtils.scala 350:94]
  assign _T_77 = 7'h11 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_78 = _T_77; // @[CFARUtils.scala 350:94]
  assign _T_81 = 7'h12 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_82 = _T_81; // @[CFARUtils.scala 350:94]
  assign _T_85 = 7'h13 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_86 = _T_85; // @[CFARUtils.scala 350:94]
  assign _T_89 = 7'h14 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_90 = _T_89; // @[CFARUtils.scala 350:94]
  assign _T_93 = 7'h15 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_94 = _T_93; // @[CFARUtils.scala 350:94]
  assign _T_97 = 7'h16 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_98 = _T_97; // @[CFARUtils.scala 350:94]
  assign _T_101 = 7'h17 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_102 = _T_101; // @[CFARUtils.scala 350:94]
  assign _T_105 = 7'h18 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_106 = _T_105; // @[CFARUtils.scala 350:94]
  assign _T_109 = 7'h19 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_110 = _T_109; // @[CFARUtils.scala 350:94]
  assign _T_113 = 7'h1a <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_114 = _T_113; // @[CFARUtils.scala 350:94]
  assign _T_117 = 7'h1b <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_118 = _T_117; // @[CFARUtils.scala 350:94]
  assign _T_121 = 7'h1c <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_122 = _T_121; // @[CFARUtils.scala 350:94]
  assign _T_125 = 7'h1d <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_126 = _T_125; // @[CFARUtils.scala 350:94]
  assign _T_129 = 7'h1e <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_130 = _T_129; // @[CFARUtils.scala 350:94]
  assign _T_133 = 7'h1f <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_134 = _T_133; // @[CFARUtils.scala 350:94]
  assign _T_137 = 7'h20 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_138 = _T_137; // @[CFARUtils.scala 350:94]
  assign _T_141 = 7'h21 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_142 = _T_141; // @[CFARUtils.scala 350:94]
  assign _T_145 = 7'h22 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_146 = _T_145; // @[CFARUtils.scala 350:94]
  assign _T_149 = 7'h23 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_150 = _T_149; // @[CFARUtils.scala 350:94]
  assign _T_153 = 7'h24 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_154 = _T_153; // @[CFARUtils.scala 350:94]
  assign _T_157 = 7'h25 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_158 = _T_157; // @[CFARUtils.scala 350:94]
  assign _T_161 = 7'h26 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_162 = _T_161; // @[CFARUtils.scala 350:94]
  assign _T_165 = 7'h27 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_166 = _T_165; // @[CFARUtils.scala 350:94]
  assign _T_169 = 7'h28 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_170 = _T_169; // @[CFARUtils.scala 350:94]
  assign _T_173 = 7'h29 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_174 = _T_173; // @[CFARUtils.scala 350:94]
  assign _T_177 = 7'h2a <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_178 = _T_177; // @[CFARUtils.scala 350:94]
  assign _T_181 = 7'h2b <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_182 = _T_181; // @[CFARUtils.scala 350:94]
  assign _T_185 = 7'h2c <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_186 = _T_185; // @[CFARUtils.scala 350:94]
  assign _T_189 = 7'h2d <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_190 = _T_189; // @[CFARUtils.scala 350:94]
  assign _T_193 = 7'h2e <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_194 = _T_193; // @[CFARUtils.scala 350:94]
  assign _T_197 = 7'h2f <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_198 = _T_197; // @[CFARUtils.scala 350:94]
  assign _T_201 = 7'h30 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_202 = _T_201; // @[CFARUtils.scala 350:94]
  assign _T_205 = 7'h31 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_206 = _T_205; // @[CFARUtils.scala 350:94]
  assign _T_209 = 7'h32 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_210 = _T_209; // @[CFARUtils.scala 350:94]
  assign _T_213 = 7'h33 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_214 = _T_213; // @[CFARUtils.scala 350:94]
  assign _T_217 = 7'h34 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_218 = _T_217; // @[CFARUtils.scala 350:94]
  assign _T_221 = 7'h35 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_222 = _T_221; // @[CFARUtils.scala 350:94]
  assign _T_225 = 7'h36 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_226 = _T_225; // @[CFARUtils.scala 350:94]
  assign _T_229 = 7'h37 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_230 = _T_229; // @[CFARUtils.scala 350:94]
  assign _T_233 = 7'h38 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_234 = _T_233; // @[CFARUtils.scala 350:94]
  assign _T_237 = 7'h39 <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_238 = _T_237; // @[CFARUtils.scala 350:94]
  assign _T_241 = 7'h3a <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_242 = _T_241; // @[CFARUtils.scala 350:94]
  assign _T_245 = 7'h3b <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_246 = _T_245; // @[CFARUtils.scala 350:94]
  assign _T_249 = 7'h3c <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_250 = _T_249; // @[CFARUtils.scala 350:94]
  assign _T_253 = 7'h3d <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_254 = _T_253; // @[CFARUtils.scala 350:94]
  assign _T_257 = 7'h3e <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_258 = _T_257; // @[CFARUtils.scala 350:94]
  assign _T_261 = 7'h3f <= _T_8; // @[CFARUtils.scala 350:78]
  assign _T_262 = _T_261; // @[CFARUtils.scala 350:94]
  assign activeRegs_63 = _T_261; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_263 = _T_262 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_62 = _T_257; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_264 = _T_258 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_61 = _T_253; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_265 = _T_254 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_60 = _T_249; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_266 = _T_250 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_59 = _T_245; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_267 = _T_246 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_58 = _T_241; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_268 = _T_242 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_57 = _T_237; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_269 = _T_238 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_56 = _T_233; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_270 = _T_234 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_55 = _T_229; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_271 = _T_230 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_54 = _T_225; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_272 = _T_226 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_53 = _T_221; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_273 = _T_222 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_52 = _T_217; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_274 = _T_218 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_51 = _T_213; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_275 = _T_214 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_50 = _T_209; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_276 = _T_210 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_49 = _T_205; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_277 = _T_206 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_48 = _T_201; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_278 = _T_202 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_47 = _T_197; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_279 = _T_198 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_46 = _T_193; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_280 = _T_194 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_45 = _T_189; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_281 = _T_190 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_44 = _T_185; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_282 = _T_186 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_43 = _T_181; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_283 = _T_182 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_42 = _T_177; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_284 = _T_178 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_41 = _T_173; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_285 = _T_174 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_40 = _T_169; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_286 = _T_170 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_39 = _T_165; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_287 = _T_166 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_38 = _T_161; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_288 = _T_162 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_37 = _T_157; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_289 = _T_158 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_36 = _T_153; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_290 = _T_154 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_35 = _T_149; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_291 = _T_150 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_34 = _T_145; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_292 = _T_146 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_33 = _T_141; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_293 = _T_142 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_32 = _T_137; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_294 = _T_138 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_31 = _T_133; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_295 = _T_134 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_30 = _T_129; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_296 = _T_130 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_29 = _T_125; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_297 = _T_126 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_28 = _T_121; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_298 = _T_122 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_27 = _T_117; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_299 = _T_118 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_26 = _T_113; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_300 = _T_114 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_25 = _T_109; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_301 = _T_110 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_24 = _T_105; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_302 = _T_106 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_23 = _T_101; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_303 = _T_102 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_22 = _T_97; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_304 = _T_98 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_21 = _T_93; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_305 = _T_94 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_20 = _T_89; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_306 = _T_90 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_19 = _T_85; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_307 = _T_86 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_18 = _T_81; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_308 = _T_82 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_17 = _T_77; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_309 = _T_78 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_16 = _T_73; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_310 = _T_74 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_15 = _T_69; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_311 = _T_70 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_14 = _T_65; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_312 = _T_66 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_13 = _T_61; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_313 = _T_62 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_12 = _T_57; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_314 = _T_58 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_11 = _T_53; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_315 = _T_54 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_10 = _T_49; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_316 = _T_50 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_9 = _T_45; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_317 = _T_46 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_8 = _T_41; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_318 = _T_42 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_7 = _T_37; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_319 = _T_38 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_6 = _T_33; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_320 = _T_34 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_5 = _T_29; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_321 = _T_30 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_4 = _T_25; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_322 = _T_26 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_3 = _T_21; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_323 = _T_22 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_2 = _T_17; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_324 = _T_18 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_1 = _T_13; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_325 = _T_14 & en; // @[CFARUtils.scala 319:37]
  assign activeRegs_0 = 1'h1; // @[CFARUtils.scala 347:26 CFARUtils.scala 350:66]
  assign _T_326 = _T_9 & en; // @[CFARUtils.scala 319:37]
  assign _T_395 = io_lastIn & _T_1; // @[CFARUtils.scala 392:19]
  assign _GEN_64 = _T_395 | last; // @[CFARUtils.scala 392:36]
  assign _T_398 = cntIn + 7'h1; // @[CFARUtils.scala 397:20]
  assign _T_399 = io_depth > 7'h1; // @[CFARUtils.scala 400:18]
  assign _T_402 = cntIn == _T_8; // @[CFARUtils.scala 401:17]
  assign _T_404 = _T_402 & _T_1; // @[CFARUtils.scala 401:36]
  assign _GEN_66 = _T_404 | InitialInDone; // @[CFARUtils.scala 401:53]
  assign _T_406 = io_depth == 7'h1; // @[CFARUtils.scala 406:36]
  assign _T_407 = _T_1 & _T_406; // @[CFARUtils.scala 406:24]
  assign _GEN_67 = _T_407 | InitialInDone; // @[CFARUtils.scala 406:45]
  assign _T_409 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_672 = _T_261 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_673 = _T_257 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_674 = _T_253 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_675 = _T_249 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_676 = _T_245 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_677 = _T_241 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_678 = _T_237 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_679 = _T_233 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_680 = _T_229 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_681 = _T_225 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_682 = _T_221 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_683 = _T_217 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_684 = _T_213 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_685 = _T_209 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_686 = _T_205 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_687 = _T_201 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_688 = _T_197 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_689 = _T_193 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_690 = _T_189 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_691 = _T_185 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_692 = _T_181 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_693 = _T_177 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_694 = _T_173 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_695 = _T_169 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_696 = _T_165 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_697 = _T_161 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_698 = _T_157 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_699 = _T_153 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_700 = _T_149 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_701 = _T_145 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_702 = _T_141 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_703 = _T_137 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_704 = _T_133 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_705 = _T_129 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_706 = _T_125 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_707 = _T_121 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_708 = _T_117 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_709 = _T_113 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_710 = _T_109 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_711 = _T_105 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_712 = _T_101 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_713 = _T_97 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_714 = _T_93 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_715 = _T_89 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_716 = _T_85 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_717 = _T_81 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_718 = _T_77 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_719 = _T_73 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_720 = _T_69 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_721 = _T_65 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_722 = _T_61 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_723 = _T_57 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_724 = _T_53 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_725 = _T_49 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_726 = _T_45 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_727 = _T_41 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_728 = _T_37 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_729 = _T_33 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_730 = _T_29 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_731 = _T_25 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_732 = _T_21 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_733 = _T_17 & _T_409; // @[CFARUtils.scala 319:37]
  assign _T_734 = _T_13 & _T_409; // @[CFARUtils.scala 319:37]
  assign _GEN_134 = 6'h1 == _T_8[5:0] ? _T_737 : _T_736; // @[CFARUtils.scala 414:17]
  assign _GEN_135 = 6'h2 == _T_8[5:0] ? _T_738 : _GEN_134; // @[CFARUtils.scala 414:17]
  assign _GEN_136 = 6'h3 == _T_8[5:0] ? _T_739 : _GEN_135; // @[CFARUtils.scala 414:17]
  assign _GEN_137 = 6'h4 == _T_8[5:0] ? _T_740 : _GEN_136; // @[CFARUtils.scala 414:17]
  assign _GEN_138 = 6'h5 == _T_8[5:0] ? _T_741 : _GEN_137; // @[CFARUtils.scala 414:17]
  assign _GEN_139 = 6'h6 == _T_8[5:0] ? _T_742 : _GEN_138; // @[CFARUtils.scala 414:17]
  assign _GEN_140 = 6'h7 == _T_8[5:0] ? _T_743 : _GEN_139; // @[CFARUtils.scala 414:17]
  assign _GEN_141 = 6'h8 == _T_8[5:0] ? _T_744 : _GEN_140; // @[CFARUtils.scala 414:17]
  assign _GEN_142 = 6'h9 == _T_8[5:0] ? _T_745 : _GEN_141; // @[CFARUtils.scala 414:17]
  assign _GEN_143 = 6'ha == _T_8[5:0] ? _T_746 : _GEN_142; // @[CFARUtils.scala 414:17]
  assign _GEN_144 = 6'hb == _T_8[5:0] ? _T_747 : _GEN_143; // @[CFARUtils.scala 414:17]
  assign _GEN_145 = 6'hc == _T_8[5:0] ? _T_748 : _GEN_144; // @[CFARUtils.scala 414:17]
  assign _GEN_146 = 6'hd == _T_8[5:0] ? _T_749 : _GEN_145; // @[CFARUtils.scala 414:17]
  assign _GEN_147 = 6'he == _T_8[5:0] ? _T_750 : _GEN_146; // @[CFARUtils.scala 414:17]
  assign _GEN_148 = 6'hf == _T_8[5:0] ? _T_751 : _GEN_147; // @[CFARUtils.scala 414:17]
  assign _GEN_149 = 6'h10 == _T_8[5:0] ? _T_752 : _GEN_148; // @[CFARUtils.scala 414:17]
  assign _GEN_150 = 6'h11 == _T_8[5:0] ? _T_753 : _GEN_149; // @[CFARUtils.scala 414:17]
  assign _GEN_151 = 6'h12 == _T_8[5:0] ? _T_754 : _GEN_150; // @[CFARUtils.scala 414:17]
  assign _GEN_152 = 6'h13 == _T_8[5:0] ? _T_755 : _GEN_151; // @[CFARUtils.scala 414:17]
  assign _GEN_153 = 6'h14 == _T_8[5:0] ? _T_756 : _GEN_152; // @[CFARUtils.scala 414:17]
  assign _GEN_154 = 6'h15 == _T_8[5:0] ? _T_757 : _GEN_153; // @[CFARUtils.scala 414:17]
  assign _GEN_155 = 6'h16 == _T_8[5:0] ? _T_758 : _GEN_154; // @[CFARUtils.scala 414:17]
  assign _GEN_156 = 6'h17 == _T_8[5:0] ? _T_759 : _GEN_155; // @[CFARUtils.scala 414:17]
  assign _GEN_157 = 6'h18 == _T_8[5:0] ? _T_760 : _GEN_156; // @[CFARUtils.scala 414:17]
  assign _GEN_158 = 6'h19 == _T_8[5:0] ? _T_761 : _GEN_157; // @[CFARUtils.scala 414:17]
  assign _GEN_159 = 6'h1a == _T_8[5:0] ? _T_762 : _GEN_158; // @[CFARUtils.scala 414:17]
  assign _GEN_160 = 6'h1b == _T_8[5:0] ? _T_763 : _GEN_159; // @[CFARUtils.scala 414:17]
  assign _GEN_161 = 6'h1c == _T_8[5:0] ? _T_764 : _GEN_160; // @[CFARUtils.scala 414:17]
  assign _GEN_162 = 6'h1d == _T_8[5:0] ? _T_765 : _GEN_161; // @[CFARUtils.scala 414:17]
  assign _GEN_163 = 6'h1e == _T_8[5:0] ? _T_766 : _GEN_162; // @[CFARUtils.scala 414:17]
  assign _GEN_164 = 6'h1f == _T_8[5:0] ? _T_767 : _GEN_163; // @[CFARUtils.scala 414:17]
  assign _GEN_165 = 6'h20 == _T_8[5:0] ? _T_768 : _GEN_164; // @[CFARUtils.scala 414:17]
  assign _GEN_166 = 6'h21 == _T_8[5:0] ? _T_769 : _GEN_165; // @[CFARUtils.scala 414:17]
  assign _GEN_167 = 6'h22 == _T_8[5:0] ? _T_770 : _GEN_166; // @[CFARUtils.scala 414:17]
  assign _GEN_168 = 6'h23 == _T_8[5:0] ? _T_771 : _GEN_167; // @[CFARUtils.scala 414:17]
  assign _GEN_169 = 6'h24 == _T_8[5:0] ? _T_772 : _GEN_168; // @[CFARUtils.scala 414:17]
  assign _GEN_170 = 6'h25 == _T_8[5:0] ? _T_773 : _GEN_169; // @[CFARUtils.scala 414:17]
  assign _GEN_171 = 6'h26 == _T_8[5:0] ? _T_774 : _GEN_170; // @[CFARUtils.scala 414:17]
  assign _GEN_172 = 6'h27 == _T_8[5:0] ? _T_775 : _GEN_171; // @[CFARUtils.scala 414:17]
  assign _GEN_173 = 6'h28 == _T_8[5:0] ? _T_776 : _GEN_172; // @[CFARUtils.scala 414:17]
  assign _GEN_174 = 6'h29 == _T_8[5:0] ? _T_777 : _GEN_173; // @[CFARUtils.scala 414:17]
  assign _GEN_175 = 6'h2a == _T_8[5:0] ? _T_778 : _GEN_174; // @[CFARUtils.scala 414:17]
  assign _GEN_176 = 6'h2b == _T_8[5:0] ? _T_779 : _GEN_175; // @[CFARUtils.scala 414:17]
  assign _GEN_177 = 6'h2c == _T_8[5:0] ? _T_780 : _GEN_176; // @[CFARUtils.scala 414:17]
  assign _GEN_178 = 6'h2d == _T_8[5:0] ? _T_781 : _GEN_177; // @[CFARUtils.scala 414:17]
  assign _GEN_179 = 6'h2e == _T_8[5:0] ? _T_782 : _GEN_178; // @[CFARUtils.scala 414:17]
  assign _GEN_180 = 6'h2f == _T_8[5:0] ? _T_783 : _GEN_179; // @[CFARUtils.scala 414:17]
  assign _GEN_181 = 6'h30 == _T_8[5:0] ? _T_784 : _GEN_180; // @[CFARUtils.scala 414:17]
  assign _GEN_182 = 6'h31 == _T_8[5:0] ? _T_785 : _GEN_181; // @[CFARUtils.scala 414:17]
  assign _GEN_183 = 6'h32 == _T_8[5:0] ? _T_786 : _GEN_182; // @[CFARUtils.scala 414:17]
  assign _GEN_184 = 6'h33 == _T_8[5:0] ? _T_787 : _GEN_183; // @[CFARUtils.scala 414:17]
  assign _GEN_185 = 6'h34 == _T_8[5:0] ? _T_788 : _GEN_184; // @[CFARUtils.scala 414:17]
  assign _GEN_186 = 6'h35 == _T_8[5:0] ? _T_789 : _GEN_185; // @[CFARUtils.scala 414:17]
  assign _GEN_187 = 6'h36 == _T_8[5:0] ? _T_790 : _GEN_186; // @[CFARUtils.scala 414:17]
  assign _GEN_188 = 6'h37 == _T_8[5:0] ? _T_791 : _GEN_187; // @[CFARUtils.scala 414:17]
  assign _GEN_189 = 6'h38 == _T_8[5:0] ? _T_792 : _GEN_188; // @[CFARUtils.scala 414:17]
  assign _GEN_190 = 6'h39 == _T_8[5:0] ? _T_793 : _GEN_189; // @[CFARUtils.scala 414:17]
  assign _GEN_191 = 6'h3a == _T_8[5:0] ? _T_794 : _GEN_190; // @[CFARUtils.scala 414:17]
  assign _GEN_192 = 6'h3b == _T_8[5:0] ? _T_795 : _GEN_191; // @[CFARUtils.scala 414:17]
  assign _GEN_193 = 6'h3c == _T_8[5:0] ? _T_796 : _GEN_192; // @[CFARUtils.scala 414:17]
  assign _GEN_194 = 6'h3d == _T_8[5:0] ? _T_797 : _GEN_193; // @[CFARUtils.scala 414:17]
  assign _GEN_195 = 6'h3e == _T_8[5:0] ? _T_798 : _GEN_194; // @[CFARUtils.scala 414:17]
  assign _GEN_196 = 6'h3f == _T_8[5:0] ? _T_799 : _GEN_195; // @[CFARUtils.scala 414:17]
  assign _T_804 = _GEN_196 & _T_409; // @[CFARUtils.scala 414:17]
  assign _T_808 = ~last; // @[CFARUtils.scala 421:36]
  assign _T_810 = io_depth == 7'h0; // @[CFARUtils.scala 429:37]
  assign _T_812 = io_out_ready & _T_808; // @[CFARUtils.scala 429:73]
  assign _T_821 = InitialInDone & io_in_valid; // @[CFARUtils.scala 436:70]
  assign _T_822 = last & en; // @[CFARUtils.scala 436:94]
  assign _T_823 = _T_821 | _T_822; // @[CFARUtils.scala 436:85]
  assign io_in_ready = _T_810 ? io_out_ready : _T_812; // @[CFARUtils.scala 429:20]
  assign io_out_valid = _T_810 ? io_in_valid : _T_823; // @[CFARUtils.scala 436:18]
  assign io_parallelOut_0 = adjShiftRegOut_0; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_1 = adjShiftRegOut_1; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_2 = adjShiftRegOut_2; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_3 = adjShiftRegOut_3; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_4 = adjShiftRegOut_4; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_5 = adjShiftRegOut_5; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_6 = adjShiftRegOut_6; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_7 = adjShiftRegOut_7; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_8 = adjShiftRegOut_8; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_9 = adjShiftRegOut_9; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_10 = adjShiftRegOut_10; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_11 = adjShiftRegOut_11; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_12 = adjShiftRegOut_12; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_13 = adjShiftRegOut_13; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_14 = adjShiftRegOut_14; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_15 = adjShiftRegOut_15; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_16 = adjShiftRegOut_16; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_17 = adjShiftRegOut_17; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_18 = adjShiftRegOut_18; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_19 = adjShiftRegOut_19; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_20 = adjShiftRegOut_20; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_21 = adjShiftRegOut_21; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_22 = adjShiftRegOut_22; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_23 = adjShiftRegOut_23; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_24 = adjShiftRegOut_24; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_25 = adjShiftRegOut_25; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_26 = adjShiftRegOut_26; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_27 = adjShiftRegOut_27; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_28 = adjShiftRegOut_28; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_29 = adjShiftRegOut_29; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_30 = adjShiftRegOut_30; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_31 = adjShiftRegOut_31; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_32 = adjShiftRegOut_32; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_33 = adjShiftRegOut_33; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_34 = adjShiftRegOut_34; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_35 = adjShiftRegOut_35; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_36 = adjShiftRegOut_36; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_37 = adjShiftRegOut_37; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_38 = adjShiftRegOut_38; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_39 = adjShiftRegOut_39; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_40 = adjShiftRegOut_40; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_41 = adjShiftRegOut_41; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_42 = adjShiftRegOut_42; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_43 = adjShiftRegOut_43; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_44 = adjShiftRegOut_44; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_45 = adjShiftRegOut_45; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_46 = adjShiftRegOut_46; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_47 = adjShiftRegOut_47; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_48 = adjShiftRegOut_48; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_49 = adjShiftRegOut_49; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_50 = adjShiftRegOut_50; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_51 = adjShiftRegOut_51; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_52 = adjShiftRegOut_52; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_53 = adjShiftRegOut_53; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_54 = adjShiftRegOut_54; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_55 = adjShiftRegOut_55; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_56 = adjShiftRegOut_56; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_57 = adjShiftRegOut_57; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_58 = adjShiftRegOut_58; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_59 = adjShiftRegOut_59; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_60 = adjShiftRegOut_60; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_61 = adjShiftRegOut_61; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_62 = adjShiftRegOut_62; // @[CFARUtils.scala 434:18]
  assign io_parallelOut_63 = adjShiftRegOut_63; // @[CFARUtils.scala 434:18]
  assign io_cnt = cntIn; // @[CFARUtils.scala 438:16]
  assign io_regFull = InitialInDone & _T_808; // @[CFARUtils.scala 421:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  InitialInDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  last = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  adjShiftRegOut_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  adjShiftRegOut_1 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  adjShiftRegOut_2 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  adjShiftRegOut_3 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  adjShiftRegOut_4 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  adjShiftRegOut_5 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  adjShiftRegOut_6 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  adjShiftRegOut_7 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  adjShiftRegOut_8 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  adjShiftRegOut_9 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  adjShiftRegOut_10 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  adjShiftRegOut_11 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  adjShiftRegOut_12 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  adjShiftRegOut_13 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  adjShiftRegOut_14 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  adjShiftRegOut_15 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  adjShiftRegOut_16 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  adjShiftRegOut_17 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  adjShiftRegOut_18 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  adjShiftRegOut_19 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  adjShiftRegOut_20 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  adjShiftRegOut_21 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  adjShiftRegOut_22 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  adjShiftRegOut_23 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  adjShiftRegOut_24 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  adjShiftRegOut_25 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  adjShiftRegOut_26 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  adjShiftRegOut_27 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  adjShiftRegOut_28 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  adjShiftRegOut_29 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  adjShiftRegOut_30 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  adjShiftRegOut_31 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  adjShiftRegOut_32 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  adjShiftRegOut_33 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  adjShiftRegOut_34 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  adjShiftRegOut_35 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  adjShiftRegOut_36 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  adjShiftRegOut_37 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  adjShiftRegOut_38 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  adjShiftRegOut_39 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  adjShiftRegOut_40 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  adjShiftRegOut_41 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  adjShiftRegOut_42 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  adjShiftRegOut_43 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  adjShiftRegOut_44 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  adjShiftRegOut_45 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  adjShiftRegOut_46 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  adjShiftRegOut_47 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  adjShiftRegOut_48 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  adjShiftRegOut_49 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  adjShiftRegOut_50 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  adjShiftRegOut_51 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  adjShiftRegOut_52 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  adjShiftRegOut_53 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  adjShiftRegOut_54 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  adjShiftRegOut_55 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  adjShiftRegOut_56 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  adjShiftRegOut_57 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  adjShiftRegOut_58 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  adjShiftRegOut_59 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  adjShiftRegOut_60 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  adjShiftRegOut_61 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  adjShiftRegOut_62 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  adjShiftRegOut_63 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  cntIn = _RAND_66[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_736 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_737 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_738 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_739 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_740 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_741 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_742 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_743 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_744 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_745 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_746 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_747 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_748 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_749 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_750 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_751 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_752 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_753 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_754 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_755 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_756 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_757 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_758 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_759 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_760 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_761 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_762 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_763 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_764 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_765 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_766 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_767 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_768 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_769 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_770 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_771 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_772 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_773 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_774 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_775 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_776 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_777 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_778 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_779 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_780 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_781 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_782 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_783 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_784 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_785 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_786 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_787 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_788 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_789 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_790 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_791 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_792 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_793 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_794 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_795 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_796 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_797 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_798 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_799 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      InitialInDone <= 1'h0;
    end else if (_T_804) begin
      InitialInDone <= 1'h0;
    end else if (_T_399) begin
      InitialInDone <= _GEN_66;
    end else begin
      InitialInDone <= _GEN_67;
    end
    if (reset) begin
      last <= 1'h0;
    end else if (_T_804) begin
      last <= 1'h0;
    end else begin
      last <= _GEN_64;
    end
    if (reset) begin
      adjShiftRegOut_0 <= 16'sh0;
    end else if (_T_326) begin
      adjShiftRegOut_0 <= io_in_bits;
    end
    if (reset) begin
      adjShiftRegOut_1 <= 16'sh0;
    end else if (_T_325) begin
      adjShiftRegOut_1 <= adjShiftRegOut_0;
    end
    if (reset) begin
      adjShiftRegOut_2 <= 16'sh0;
    end else if (_T_324) begin
      adjShiftRegOut_2 <= adjShiftRegOut_1;
    end
    if (reset) begin
      adjShiftRegOut_3 <= 16'sh0;
    end else if (_T_323) begin
      adjShiftRegOut_3 <= adjShiftRegOut_2;
    end
    if (reset) begin
      adjShiftRegOut_4 <= 16'sh0;
    end else if (_T_322) begin
      adjShiftRegOut_4 <= adjShiftRegOut_3;
    end
    if (reset) begin
      adjShiftRegOut_5 <= 16'sh0;
    end else if (_T_321) begin
      adjShiftRegOut_5 <= adjShiftRegOut_4;
    end
    if (reset) begin
      adjShiftRegOut_6 <= 16'sh0;
    end else if (_T_320) begin
      adjShiftRegOut_6 <= adjShiftRegOut_5;
    end
    if (reset) begin
      adjShiftRegOut_7 <= 16'sh0;
    end else if (_T_319) begin
      adjShiftRegOut_7 <= adjShiftRegOut_6;
    end
    if (reset) begin
      adjShiftRegOut_8 <= 16'sh0;
    end else if (_T_318) begin
      adjShiftRegOut_8 <= adjShiftRegOut_7;
    end
    if (reset) begin
      adjShiftRegOut_9 <= 16'sh0;
    end else if (_T_317) begin
      adjShiftRegOut_9 <= adjShiftRegOut_8;
    end
    if (reset) begin
      adjShiftRegOut_10 <= 16'sh0;
    end else if (_T_316) begin
      adjShiftRegOut_10 <= adjShiftRegOut_9;
    end
    if (reset) begin
      adjShiftRegOut_11 <= 16'sh0;
    end else if (_T_315) begin
      adjShiftRegOut_11 <= adjShiftRegOut_10;
    end
    if (reset) begin
      adjShiftRegOut_12 <= 16'sh0;
    end else if (_T_314) begin
      adjShiftRegOut_12 <= adjShiftRegOut_11;
    end
    if (reset) begin
      adjShiftRegOut_13 <= 16'sh0;
    end else if (_T_313) begin
      adjShiftRegOut_13 <= adjShiftRegOut_12;
    end
    if (reset) begin
      adjShiftRegOut_14 <= 16'sh0;
    end else if (_T_312) begin
      adjShiftRegOut_14 <= adjShiftRegOut_13;
    end
    if (reset) begin
      adjShiftRegOut_15 <= 16'sh0;
    end else if (_T_311) begin
      adjShiftRegOut_15 <= adjShiftRegOut_14;
    end
    if (reset) begin
      adjShiftRegOut_16 <= 16'sh0;
    end else if (_T_310) begin
      adjShiftRegOut_16 <= adjShiftRegOut_15;
    end
    if (reset) begin
      adjShiftRegOut_17 <= 16'sh0;
    end else if (_T_309) begin
      adjShiftRegOut_17 <= adjShiftRegOut_16;
    end
    if (reset) begin
      adjShiftRegOut_18 <= 16'sh0;
    end else if (_T_308) begin
      adjShiftRegOut_18 <= adjShiftRegOut_17;
    end
    if (reset) begin
      adjShiftRegOut_19 <= 16'sh0;
    end else if (_T_307) begin
      adjShiftRegOut_19 <= adjShiftRegOut_18;
    end
    if (reset) begin
      adjShiftRegOut_20 <= 16'sh0;
    end else if (_T_306) begin
      adjShiftRegOut_20 <= adjShiftRegOut_19;
    end
    if (reset) begin
      adjShiftRegOut_21 <= 16'sh0;
    end else if (_T_305) begin
      adjShiftRegOut_21 <= adjShiftRegOut_20;
    end
    if (reset) begin
      adjShiftRegOut_22 <= 16'sh0;
    end else if (_T_304) begin
      adjShiftRegOut_22 <= adjShiftRegOut_21;
    end
    if (reset) begin
      adjShiftRegOut_23 <= 16'sh0;
    end else if (_T_303) begin
      adjShiftRegOut_23 <= adjShiftRegOut_22;
    end
    if (reset) begin
      adjShiftRegOut_24 <= 16'sh0;
    end else if (_T_302) begin
      adjShiftRegOut_24 <= adjShiftRegOut_23;
    end
    if (reset) begin
      adjShiftRegOut_25 <= 16'sh0;
    end else if (_T_301) begin
      adjShiftRegOut_25 <= adjShiftRegOut_24;
    end
    if (reset) begin
      adjShiftRegOut_26 <= 16'sh0;
    end else if (_T_300) begin
      adjShiftRegOut_26 <= adjShiftRegOut_25;
    end
    if (reset) begin
      adjShiftRegOut_27 <= 16'sh0;
    end else if (_T_299) begin
      adjShiftRegOut_27 <= adjShiftRegOut_26;
    end
    if (reset) begin
      adjShiftRegOut_28 <= 16'sh0;
    end else if (_T_298) begin
      adjShiftRegOut_28 <= adjShiftRegOut_27;
    end
    if (reset) begin
      adjShiftRegOut_29 <= 16'sh0;
    end else if (_T_297) begin
      adjShiftRegOut_29 <= adjShiftRegOut_28;
    end
    if (reset) begin
      adjShiftRegOut_30 <= 16'sh0;
    end else if (_T_296) begin
      adjShiftRegOut_30 <= adjShiftRegOut_29;
    end
    if (reset) begin
      adjShiftRegOut_31 <= 16'sh0;
    end else if (_T_295) begin
      adjShiftRegOut_31 <= adjShiftRegOut_30;
    end
    if (reset) begin
      adjShiftRegOut_32 <= 16'sh0;
    end else if (_T_294) begin
      adjShiftRegOut_32 <= adjShiftRegOut_31;
    end
    if (reset) begin
      adjShiftRegOut_33 <= 16'sh0;
    end else if (_T_293) begin
      adjShiftRegOut_33 <= adjShiftRegOut_32;
    end
    if (reset) begin
      adjShiftRegOut_34 <= 16'sh0;
    end else if (_T_292) begin
      adjShiftRegOut_34 <= adjShiftRegOut_33;
    end
    if (reset) begin
      adjShiftRegOut_35 <= 16'sh0;
    end else if (_T_291) begin
      adjShiftRegOut_35 <= adjShiftRegOut_34;
    end
    if (reset) begin
      adjShiftRegOut_36 <= 16'sh0;
    end else if (_T_290) begin
      adjShiftRegOut_36 <= adjShiftRegOut_35;
    end
    if (reset) begin
      adjShiftRegOut_37 <= 16'sh0;
    end else if (_T_289) begin
      adjShiftRegOut_37 <= adjShiftRegOut_36;
    end
    if (reset) begin
      adjShiftRegOut_38 <= 16'sh0;
    end else if (_T_288) begin
      adjShiftRegOut_38 <= adjShiftRegOut_37;
    end
    if (reset) begin
      adjShiftRegOut_39 <= 16'sh0;
    end else if (_T_287) begin
      adjShiftRegOut_39 <= adjShiftRegOut_38;
    end
    if (reset) begin
      adjShiftRegOut_40 <= 16'sh0;
    end else if (_T_286) begin
      adjShiftRegOut_40 <= adjShiftRegOut_39;
    end
    if (reset) begin
      adjShiftRegOut_41 <= 16'sh0;
    end else if (_T_285) begin
      adjShiftRegOut_41 <= adjShiftRegOut_40;
    end
    if (reset) begin
      adjShiftRegOut_42 <= 16'sh0;
    end else if (_T_284) begin
      adjShiftRegOut_42 <= adjShiftRegOut_41;
    end
    if (reset) begin
      adjShiftRegOut_43 <= 16'sh0;
    end else if (_T_283) begin
      adjShiftRegOut_43 <= adjShiftRegOut_42;
    end
    if (reset) begin
      adjShiftRegOut_44 <= 16'sh0;
    end else if (_T_282) begin
      adjShiftRegOut_44 <= adjShiftRegOut_43;
    end
    if (reset) begin
      adjShiftRegOut_45 <= 16'sh0;
    end else if (_T_281) begin
      adjShiftRegOut_45 <= adjShiftRegOut_44;
    end
    if (reset) begin
      adjShiftRegOut_46 <= 16'sh0;
    end else if (_T_280) begin
      adjShiftRegOut_46 <= adjShiftRegOut_45;
    end
    if (reset) begin
      adjShiftRegOut_47 <= 16'sh0;
    end else if (_T_279) begin
      adjShiftRegOut_47 <= adjShiftRegOut_46;
    end
    if (reset) begin
      adjShiftRegOut_48 <= 16'sh0;
    end else if (_T_278) begin
      adjShiftRegOut_48 <= adjShiftRegOut_47;
    end
    if (reset) begin
      adjShiftRegOut_49 <= 16'sh0;
    end else if (_T_277) begin
      adjShiftRegOut_49 <= adjShiftRegOut_48;
    end
    if (reset) begin
      adjShiftRegOut_50 <= 16'sh0;
    end else if (_T_276) begin
      adjShiftRegOut_50 <= adjShiftRegOut_49;
    end
    if (reset) begin
      adjShiftRegOut_51 <= 16'sh0;
    end else if (_T_275) begin
      adjShiftRegOut_51 <= adjShiftRegOut_50;
    end
    if (reset) begin
      adjShiftRegOut_52 <= 16'sh0;
    end else if (_T_274) begin
      adjShiftRegOut_52 <= adjShiftRegOut_51;
    end
    if (reset) begin
      adjShiftRegOut_53 <= 16'sh0;
    end else if (_T_273) begin
      adjShiftRegOut_53 <= adjShiftRegOut_52;
    end
    if (reset) begin
      adjShiftRegOut_54 <= 16'sh0;
    end else if (_T_272) begin
      adjShiftRegOut_54 <= adjShiftRegOut_53;
    end
    if (reset) begin
      adjShiftRegOut_55 <= 16'sh0;
    end else if (_T_271) begin
      adjShiftRegOut_55 <= adjShiftRegOut_54;
    end
    if (reset) begin
      adjShiftRegOut_56 <= 16'sh0;
    end else if (_T_270) begin
      adjShiftRegOut_56 <= adjShiftRegOut_55;
    end
    if (reset) begin
      adjShiftRegOut_57 <= 16'sh0;
    end else if (_T_269) begin
      adjShiftRegOut_57 <= adjShiftRegOut_56;
    end
    if (reset) begin
      adjShiftRegOut_58 <= 16'sh0;
    end else if (_T_268) begin
      adjShiftRegOut_58 <= adjShiftRegOut_57;
    end
    if (reset) begin
      adjShiftRegOut_59 <= 16'sh0;
    end else if (_T_267) begin
      adjShiftRegOut_59 <= adjShiftRegOut_58;
    end
    if (reset) begin
      adjShiftRegOut_60 <= 16'sh0;
    end else if (_T_266) begin
      adjShiftRegOut_60 <= adjShiftRegOut_59;
    end
    if (reset) begin
      adjShiftRegOut_61 <= 16'sh0;
    end else if (_T_265) begin
      adjShiftRegOut_61 <= adjShiftRegOut_60;
    end
    if (reset) begin
      adjShiftRegOut_62 <= 16'sh0;
    end else if (_T_264) begin
      adjShiftRegOut_62 <= adjShiftRegOut_61;
    end
    if (reset) begin
      adjShiftRegOut_63 <= 16'sh0;
    end else if (_T_263) begin
      adjShiftRegOut_63 <= adjShiftRegOut_62;
    end
    if (reset) begin
      cntIn <= 7'h0;
    end else if (_T_804) begin
      cntIn <= 7'h0;
    end else if (_T_1) begin
      cntIn <= _T_398;
    end
    if (reset) begin
      _T_736 <= 1'h0;
    end else if (_T_409) begin
      _T_736 <= _T_395;
    end
    if (reset) begin
      _T_737 <= 1'h0;
    end else if (_T_734) begin
      _T_737 <= _T_736;
    end
    if (reset) begin
      _T_738 <= 1'h0;
    end else if (_T_733) begin
      _T_738 <= _T_737;
    end
    if (reset) begin
      _T_739 <= 1'h0;
    end else if (_T_732) begin
      _T_739 <= _T_738;
    end
    if (reset) begin
      _T_740 <= 1'h0;
    end else if (_T_731) begin
      _T_740 <= _T_739;
    end
    if (reset) begin
      _T_741 <= 1'h0;
    end else if (_T_730) begin
      _T_741 <= _T_740;
    end
    if (reset) begin
      _T_742 <= 1'h0;
    end else if (_T_729) begin
      _T_742 <= _T_741;
    end
    if (reset) begin
      _T_743 <= 1'h0;
    end else if (_T_728) begin
      _T_743 <= _T_742;
    end
    if (reset) begin
      _T_744 <= 1'h0;
    end else if (_T_727) begin
      _T_744 <= _T_743;
    end
    if (reset) begin
      _T_745 <= 1'h0;
    end else if (_T_726) begin
      _T_745 <= _T_744;
    end
    if (reset) begin
      _T_746 <= 1'h0;
    end else if (_T_725) begin
      _T_746 <= _T_745;
    end
    if (reset) begin
      _T_747 <= 1'h0;
    end else if (_T_724) begin
      _T_747 <= _T_746;
    end
    if (reset) begin
      _T_748 <= 1'h0;
    end else if (_T_723) begin
      _T_748 <= _T_747;
    end
    if (reset) begin
      _T_749 <= 1'h0;
    end else if (_T_722) begin
      _T_749 <= _T_748;
    end
    if (reset) begin
      _T_750 <= 1'h0;
    end else if (_T_721) begin
      _T_750 <= _T_749;
    end
    if (reset) begin
      _T_751 <= 1'h0;
    end else if (_T_720) begin
      _T_751 <= _T_750;
    end
    if (reset) begin
      _T_752 <= 1'h0;
    end else if (_T_719) begin
      _T_752 <= _T_751;
    end
    if (reset) begin
      _T_753 <= 1'h0;
    end else if (_T_718) begin
      _T_753 <= _T_752;
    end
    if (reset) begin
      _T_754 <= 1'h0;
    end else if (_T_717) begin
      _T_754 <= _T_753;
    end
    if (reset) begin
      _T_755 <= 1'h0;
    end else if (_T_716) begin
      _T_755 <= _T_754;
    end
    if (reset) begin
      _T_756 <= 1'h0;
    end else if (_T_715) begin
      _T_756 <= _T_755;
    end
    if (reset) begin
      _T_757 <= 1'h0;
    end else if (_T_714) begin
      _T_757 <= _T_756;
    end
    if (reset) begin
      _T_758 <= 1'h0;
    end else if (_T_713) begin
      _T_758 <= _T_757;
    end
    if (reset) begin
      _T_759 <= 1'h0;
    end else if (_T_712) begin
      _T_759 <= _T_758;
    end
    if (reset) begin
      _T_760 <= 1'h0;
    end else if (_T_711) begin
      _T_760 <= _T_759;
    end
    if (reset) begin
      _T_761 <= 1'h0;
    end else if (_T_710) begin
      _T_761 <= _T_760;
    end
    if (reset) begin
      _T_762 <= 1'h0;
    end else if (_T_709) begin
      _T_762 <= _T_761;
    end
    if (reset) begin
      _T_763 <= 1'h0;
    end else if (_T_708) begin
      _T_763 <= _T_762;
    end
    if (reset) begin
      _T_764 <= 1'h0;
    end else if (_T_707) begin
      _T_764 <= _T_763;
    end
    if (reset) begin
      _T_765 <= 1'h0;
    end else if (_T_706) begin
      _T_765 <= _T_764;
    end
    if (reset) begin
      _T_766 <= 1'h0;
    end else if (_T_705) begin
      _T_766 <= _T_765;
    end
    if (reset) begin
      _T_767 <= 1'h0;
    end else if (_T_704) begin
      _T_767 <= _T_766;
    end
    if (reset) begin
      _T_768 <= 1'h0;
    end else if (_T_703) begin
      _T_768 <= _T_767;
    end
    if (reset) begin
      _T_769 <= 1'h0;
    end else if (_T_702) begin
      _T_769 <= _T_768;
    end
    if (reset) begin
      _T_770 <= 1'h0;
    end else if (_T_701) begin
      _T_770 <= _T_769;
    end
    if (reset) begin
      _T_771 <= 1'h0;
    end else if (_T_700) begin
      _T_771 <= _T_770;
    end
    if (reset) begin
      _T_772 <= 1'h0;
    end else if (_T_699) begin
      _T_772 <= _T_771;
    end
    if (reset) begin
      _T_773 <= 1'h0;
    end else if (_T_698) begin
      _T_773 <= _T_772;
    end
    if (reset) begin
      _T_774 <= 1'h0;
    end else if (_T_697) begin
      _T_774 <= _T_773;
    end
    if (reset) begin
      _T_775 <= 1'h0;
    end else if (_T_696) begin
      _T_775 <= _T_774;
    end
    if (reset) begin
      _T_776 <= 1'h0;
    end else if (_T_695) begin
      _T_776 <= _T_775;
    end
    if (reset) begin
      _T_777 <= 1'h0;
    end else if (_T_694) begin
      _T_777 <= _T_776;
    end
    if (reset) begin
      _T_778 <= 1'h0;
    end else if (_T_693) begin
      _T_778 <= _T_777;
    end
    if (reset) begin
      _T_779 <= 1'h0;
    end else if (_T_692) begin
      _T_779 <= _T_778;
    end
    if (reset) begin
      _T_780 <= 1'h0;
    end else if (_T_691) begin
      _T_780 <= _T_779;
    end
    if (reset) begin
      _T_781 <= 1'h0;
    end else if (_T_690) begin
      _T_781 <= _T_780;
    end
    if (reset) begin
      _T_782 <= 1'h0;
    end else if (_T_689) begin
      _T_782 <= _T_781;
    end
    if (reset) begin
      _T_783 <= 1'h0;
    end else if (_T_688) begin
      _T_783 <= _T_782;
    end
    if (reset) begin
      _T_784 <= 1'h0;
    end else if (_T_687) begin
      _T_784 <= _T_783;
    end
    if (reset) begin
      _T_785 <= 1'h0;
    end else if (_T_686) begin
      _T_785 <= _T_784;
    end
    if (reset) begin
      _T_786 <= 1'h0;
    end else if (_T_685) begin
      _T_786 <= _T_785;
    end
    if (reset) begin
      _T_787 <= 1'h0;
    end else if (_T_684) begin
      _T_787 <= _T_786;
    end
    if (reset) begin
      _T_788 <= 1'h0;
    end else if (_T_683) begin
      _T_788 <= _T_787;
    end
    if (reset) begin
      _T_789 <= 1'h0;
    end else if (_T_682) begin
      _T_789 <= _T_788;
    end
    if (reset) begin
      _T_790 <= 1'h0;
    end else if (_T_681) begin
      _T_790 <= _T_789;
    end
    if (reset) begin
      _T_791 <= 1'h0;
    end else if (_T_680) begin
      _T_791 <= _T_790;
    end
    if (reset) begin
      _T_792 <= 1'h0;
    end else if (_T_679) begin
      _T_792 <= _T_791;
    end
    if (reset) begin
      _T_793 <= 1'h0;
    end else if (_T_678) begin
      _T_793 <= _T_792;
    end
    if (reset) begin
      _T_794 <= 1'h0;
    end else if (_T_677) begin
      _T_794 <= _T_793;
    end
    if (reset) begin
      _T_795 <= 1'h0;
    end else if (_T_676) begin
      _T_795 <= _T_794;
    end
    if (reset) begin
      _T_796 <= 1'h0;
    end else if (_T_675) begin
      _T_796 <= _T_795;
    end
    if (reset) begin
      _T_797 <= 1'h0;
    end else if (_T_674) begin
      _T_797 <= _T_796;
    end
    if (reset) begin
      _T_798 <= 1'h0;
    end else if (_T_673) begin
      _T_798 <= _T_797;
    end
    if (reset) begin
      _T_799 <= 1'h0;
    end else if (_T_672) begin
      _T_799 <= _T_798;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:345 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 345:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[CFARUtils.scala 345:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CFARUtils.scala:330 assert(depth <= maxDepth.U)\n"); // @[CFARUtils.scala 330:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[CFARUtils.scala 330:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MinimumCircuit(
  input         clock,
  input  [19:0] io_in_0,
  input  [19:0] io_in_1,
  input  [19:0] io_in_2,
  input  [19:0] io_in_3,
  input  [19:0] io_in_4,
  input  [19:0] io_in_5,
  input  [19:0] io_in_6,
  input  [19:0] io_in_7,
  input  [19:0] io_in_8,
  input  [19:0] io_in_9,
  input  [19:0] io_in_10,
  input  [19:0] io_in_11,
  input  [19:0] io_in_12,
  input  [19:0] io_in_13,
  input  [19:0] io_in_14,
  input  [19:0] io_in_15,
  input  [4:0]  io_inSize,
  output [19:0] io_out
);
  wire  _T; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_1; // @[MinimumCircuit.scala 52:54]
  wire  _T_2; // @[MinimumCircuit.scala 28:23]
  wire  _T_3; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_4; // @[MinimumCircuit.scala 52:54]
  wire  _T_5; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_6; // @[MinimumCircuit.scala 52:54]
  wire  _T_7; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_8; // @[MinimumCircuit.scala 52:54]
  wire  _T_9; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_10; // @[MinimumCircuit.scala 52:54]
  wire  _T_11; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_12; // @[MinimumCircuit.scala 52:54]
  wire  _T_13; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_14; // @[MinimumCircuit.scala 52:54]
  wire  _T_15; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_16; // @[MinimumCircuit.scala 52:54]
  wire [19:0] _T_17; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_18; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_19; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_20; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_21; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_22; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_23; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_24; // @[MinimumCircuit.scala 30:62]
  wire  _T_25; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_26; // @[MinimumCircuit.scala 31:57]
  wire  _T_27; // @[MinimumCircuit.scala 28:23]
  wire  _T_28; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_29; // @[MinimumCircuit.scala 31:57]
  wire  _T_30; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_31; // @[MinimumCircuit.scala 31:57]
  wire  _T_32; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_33; // @[MinimumCircuit.scala 31:57]
  wire [19:0] _T_34; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_35; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_36; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_37; // @[MinimumCircuit.scala 30:62]
  wire  _T_38; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_39; // @[MinimumCircuit.scala 31:57]
  wire  _T_40; // @[MinimumCircuit.scala 28:23]
  wire  _T_41; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] _T_42; // @[MinimumCircuit.scala 31:57]
  wire [19:0] _T_43; // @[MinimumCircuit.scala 30:62]
  wire [19:0] _T_44; // @[MinimumCircuit.scala 30:62]
  wire  _T_45; // @[FixedPointTypeClass.scala 53:59]
  reg [19:0] _T_47; // @[MinimumCircuit.scala 53:41]
  reg [31:0] _RAND_0;
  wire  _T_48; // @[MinimumCircuit.scala 55:27]
  reg [19:0] _T_49; // @[MinimumCircuit.scala 57:28]
  reg [31:0] _RAND_1;
  assign _T = $signed(io_in_0) < $signed(io_in_1); // @[FixedPointTypeClass.scala 53:59]
  assign _T_1 = _T ? $signed(io_in_0) : $signed(io_in_1); // @[MinimumCircuit.scala 52:54]
  assign _T_2 = 5'h8 == io_inSize; // @[MinimumCircuit.scala 28:23]
  assign _T_3 = $signed(io_in_2) < $signed(io_in_3); // @[FixedPointTypeClass.scala 53:59]
  assign _T_4 = _T_3 ? $signed(io_in_2) : $signed(io_in_3); // @[MinimumCircuit.scala 52:54]
  assign _T_5 = $signed(io_in_4) < $signed(io_in_5); // @[FixedPointTypeClass.scala 53:59]
  assign _T_6 = _T_5 ? $signed(io_in_4) : $signed(io_in_5); // @[MinimumCircuit.scala 52:54]
  assign _T_7 = $signed(io_in_6) < $signed(io_in_7); // @[FixedPointTypeClass.scala 53:59]
  assign _T_8 = _T_7 ? $signed(io_in_6) : $signed(io_in_7); // @[MinimumCircuit.scala 52:54]
  assign _T_9 = $signed(io_in_8) < $signed(io_in_9); // @[FixedPointTypeClass.scala 53:59]
  assign _T_10 = _T_9 ? $signed(io_in_8) : $signed(io_in_9); // @[MinimumCircuit.scala 52:54]
  assign _T_11 = $signed(io_in_10) < $signed(io_in_11); // @[FixedPointTypeClass.scala 53:59]
  assign _T_12 = _T_11 ? $signed(io_in_10) : $signed(io_in_11); // @[MinimumCircuit.scala 52:54]
  assign _T_13 = $signed(io_in_12) < $signed(io_in_13); // @[FixedPointTypeClass.scala 53:59]
  assign _T_14 = _T_13 ? $signed(io_in_12) : $signed(io_in_13); // @[MinimumCircuit.scala 52:54]
  assign _T_15 = $signed(io_in_14) < $signed(io_in_15); // @[FixedPointTypeClass.scala 53:59]
  assign _T_16 = _T_15 ? $signed(io_in_14) : $signed(io_in_15); // @[MinimumCircuit.scala 52:54]
  assign _T_17 = _T_2 ? $signed(io_in_0) : $signed(_T_1); // @[MinimumCircuit.scala 30:62]
  assign _T_18 = _T_2 ? $signed(io_in_1) : $signed(_T_4); // @[MinimumCircuit.scala 30:62]
  assign _T_19 = _T_2 ? $signed(io_in_2) : $signed(_T_6); // @[MinimumCircuit.scala 30:62]
  assign _T_20 = _T_2 ? $signed(io_in_3) : $signed(_T_8); // @[MinimumCircuit.scala 30:62]
  assign _T_21 = _T_2 ? $signed(io_in_4) : $signed(_T_10); // @[MinimumCircuit.scala 30:62]
  assign _T_22 = _T_2 ? $signed(io_in_5) : $signed(_T_12); // @[MinimumCircuit.scala 30:62]
  assign _T_23 = _T_2 ? $signed(io_in_6) : $signed(_T_14); // @[MinimumCircuit.scala 30:62]
  assign _T_24 = _T_2 ? $signed(io_in_7) : $signed(_T_16); // @[MinimumCircuit.scala 30:62]
  assign _T_25 = $signed(_T_17) < $signed(_T_18); // @[FixedPointTypeClass.scala 53:59]
  assign _T_26 = _T_25 ? $signed(_T_17) : $signed(_T_18); // @[MinimumCircuit.scala 31:57]
  assign _T_27 = 5'h4 == io_inSize; // @[MinimumCircuit.scala 28:23]
  assign _T_28 = $signed(_T_19) < $signed(_T_20); // @[FixedPointTypeClass.scala 53:59]
  assign _T_29 = _T_28 ? $signed(_T_19) : $signed(_T_20); // @[MinimumCircuit.scala 31:57]
  assign _T_30 = $signed(_T_21) < $signed(_T_22); // @[FixedPointTypeClass.scala 53:59]
  assign _T_31 = _T_30 ? $signed(_T_21) : $signed(_T_22); // @[MinimumCircuit.scala 31:57]
  assign _T_32 = $signed(_T_23) < $signed(_T_24); // @[FixedPointTypeClass.scala 53:59]
  assign _T_33 = _T_32 ? $signed(_T_23) : $signed(_T_24); // @[MinimumCircuit.scala 31:57]
  assign _T_34 = _T_27 ? $signed(io_in_0) : $signed(_T_26); // @[MinimumCircuit.scala 30:62]
  assign _T_35 = _T_27 ? $signed(io_in_1) : $signed(_T_29); // @[MinimumCircuit.scala 30:62]
  assign _T_36 = _T_27 ? $signed(io_in_2) : $signed(_T_31); // @[MinimumCircuit.scala 30:62]
  assign _T_37 = _T_27 ? $signed(io_in_3) : $signed(_T_33); // @[MinimumCircuit.scala 30:62]
  assign _T_38 = $signed(_T_34) < $signed(_T_35); // @[FixedPointTypeClass.scala 53:59]
  assign _T_39 = _T_38 ? $signed(_T_34) : $signed(_T_35); // @[MinimumCircuit.scala 31:57]
  assign _T_40 = 5'h2 == io_inSize; // @[MinimumCircuit.scala 28:23]
  assign _T_41 = $signed(_T_36) < $signed(_T_37); // @[FixedPointTypeClass.scala 53:59]
  assign _T_42 = _T_41 ? $signed(_T_36) : $signed(_T_37); // @[MinimumCircuit.scala 31:57]
  assign _T_43 = _T_40 ? $signed(io_in_0) : $signed(_T_39); // @[MinimumCircuit.scala 30:62]
  assign _T_44 = _T_40 ? $signed(io_in_1) : $signed(_T_42); // @[MinimumCircuit.scala 30:62]
  assign _T_45 = $signed(_T_43) < $signed(_T_44); // @[FixedPointTypeClass.scala 53:59]
  assign _T_48 = io_inSize == 5'h1; // @[MinimumCircuit.scala 55:27]
  assign io_out = _T_48 ? $signed(_T_49) : $signed(_T_47); // @[MinimumCircuit.scala 57:18 MinimumCircuit.scala 62:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_47 = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_49 = _RAND_1[19:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_45) begin
      if (_T_40) begin
        _T_47 <= io_in_0;
      end else if (_T_38) begin
        if (_T_27) begin
          _T_47 <= io_in_0;
        end else if (_T_25) begin
          if (_T_2) begin
            _T_47 <= io_in_0;
          end else if (_T) begin
            _T_47 <= io_in_0;
          end else begin
            _T_47 <= io_in_1;
          end
        end else if (_T_2) begin
          _T_47 <= io_in_1;
        end else if (_T_3) begin
          _T_47 <= io_in_2;
        end else begin
          _T_47 <= io_in_3;
        end
      end else if (_T_27) begin
        _T_47 <= io_in_1;
      end else if (_T_28) begin
        if (_T_2) begin
          _T_47 <= io_in_2;
        end else if (_T_5) begin
          _T_47 <= io_in_4;
        end else begin
          _T_47 <= io_in_5;
        end
      end else if (_T_2) begin
        _T_47 <= io_in_3;
      end else if (_T_7) begin
        _T_47 <= io_in_6;
      end else begin
        _T_47 <= io_in_7;
      end
    end else if (_T_40) begin
      _T_47 <= io_in_1;
    end else if (_T_41) begin
      if (_T_27) begin
        _T_47 <= io_in_2;
      end else if (_T_30) begin
        if (_T_2) begin
          _T_47 <= io_in_4;
        end else if (_T_9) begin
          _T_47 <= io_in_8;
        end else begin
          _T_47 <= io_in_9;
        end
      end else if (_T_2) begin
        _T_47 <= io_in_5;
      end else if (_T_11) begin
        _T_47 <= io_in_10;
      end else begin
        _T_47 <= io_in_11;
      end
    end else if (_T_27) begin
      _T_47 <= io_in_3;
    end else if (_T_32) begin
      if (_T_2) begin
        _T_47 <= io_in_6;
      end else if (_T_13) begin
        _T_47 <= io_in_12;
      end else begin
        _T_47 <= io_in_13;
      end
    end else if (_T_2) begin
      _T_47 <= io_in_7;
    end else if (_T_15) begin
      _T_47 <= io_in_14;
    end else begin
      _T_47 <= io_in_15;
    end
    _T_49 <= io_in_0;
  end
endmodule
module Queue_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_peak,
  input  [15:0] io_enq_bits_cut,
  input  [15:0] io_enq_bits_threshold,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_peak,
  output [15:0] io_deq_bits_cut,
  output [15:0] io_deq_bits_threshold
);
  reg  _T_peak [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_peak__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_peak__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_peak__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_peak__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_peak__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_peak__T_10_en; // @[Decoupled.scala 209:24]
  reg [15:0] _T_cut [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T_cut__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_cut__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] _T_cut__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_cut__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_cut__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_cut__T_10_en; // @[Decoupled.scala 209:24]
  reg [15:0] _T_threshold [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T_threshold__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_threshold__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] _T_threshold__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_threshold__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_threshold__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_threshold__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_5;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _GEN_11; // @[Decoupled.scala 240:27]
  wire  _GEN_16; // @[Decoupled.scala 237:18]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _GEN_15; // @[Decoupled.scala 237:18]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire  _T_16; // @[Decoupled.scala 231:19]
  assign _T_peak__T_18_addr = value_1;
  assign _T_peak__T_18_data = _T_peak[_T_peak__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_peak__T_10_data = io_enq_bits_peak;
  assign _T_peak__T_10_addr = value;
  assign _T_peak__T_10_mask = 1'h1;
  assign _T_peak__T_10_en = _T_4 ? _GEN_11 : _T_6;
  assign _T_cut__T_18_addr = value_1;
  assign _T_cut__T_18_data = _T_cut[_T_cut__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_cut__T_10_data = io_enq_bits_cut;
  assign _T_cut__T_10_addr = value;
  assign _T_cut__T_10_mask = 1'h1;
  assign _T_cut__T_10_en = _T_4 ? _GEN_11 : _T_6;
  assign _T_threshold__T_18_addr = value_1;
  assign _T_threshold__T_18_data = _T_threshold[_T_threshold__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_threshold__T_10_data = io_enq_bits_threshold;
  assign _T_threshold__T_10_addr = value;
  assign _T_threshold__T_10_mask = 1'h1;
  assign _T_threshold__T_10_en = _T_4 ? _GEN_11 : _T_6;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_11 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_16 = _T_4 ? _GEN_11 : _T_6; // @[Decoupled.scala 237:18]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_15 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_15 = _GEN_16 != _GEN_15; // @[Decoupled.scala 227:16]
  assign _T_16 = ~_T_4; // @[Decoupled.scala 231:19]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_peak = _T_4 ? io_enq_bits_peak : _T_peak__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_cut = _T_4 ? $signed(io_enq_bits_cut) : $signed(_T_cut__T_18_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_threshold = _T_4 ? $signed(io_enq_bits_threshold) : $signed(_T_threshold__T_18_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_peak[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_cut[initvar] = _RAND_1[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_threshold[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_peak__T_10_en & _T_peak__T_10_mask) begin
      _T_peak[_T_peak__T_10_addr] <= _T_peak__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_cut__T_10_en & _T_cut__T_10_mask) begin
      _T_cut[_T_cut__T_10_addr] <= _T_cut__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_threshold__T_10_en & _T_threshold__T_10_mask) begin
      _T_threshold[_T_threshold__T_10_addr] <= _T_threshold__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_16) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_15) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module Queue_6(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
  reg  _T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _GEN_9; // @[Decoupled.scala 240:27]
  wire  _GEN_12; // @[Decoupled.scala 237:18]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _GEN_11; // @[Decoupled.scala 237:18]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire  _T_16; // @[Decoupled.scala 231:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = _T_4 ? _GEN_9 : _T_6;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_12 = _T_4 ? _GEN_9 : _T_6; // @[Decoupled.scala 237:18]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_11 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_15 = _GEN_12 != _GEN_11; // @[Decoupled.scala 227:16]
  assign _T_16 = ~_T_4; // @[Decoupled.scala 231:19]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = _T_4 ? io_enq_bits : _T__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_12) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_11) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module CFARCoreWithASR(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input  [9:0]  io_fftWin,
  input  [15:0] io_thresholdScaler,
  input  [2:0]  io_divSum,
  input         io_peakGrouping,
  input  [1:0]  io_cfarMode,
  input  [6:0]  io_windowCells,
  input  [3:0]  io_guardCells,
  input  [6:0]  io_subCells,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_peak,
  output [15:0] io_out_bits_cut,
  output [15:0] io_out_bits_threshold,
  output        io_lastOut,
  output [8:0]  io_fftBin
);
  wire  laggWindow_clock; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_reset; // @[CFARCoreWithASR.scala 43:30]
  wire [6:0] laggWindow_io_depth; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_io_in_ready; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_io_in_valid; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_in_bits; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_io_lastIn; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_io_out_ready; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_io_out_valid; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_out_bits; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_io_lastOut; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_0; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_1; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_2; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_3; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_4; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_5; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_6; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_7; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_8; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_9; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_10; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_11; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_12; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_13; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_14; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_15; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_16; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_17; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_18; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_19; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_20; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_21; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_22; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_23; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_24; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_25; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_26; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_27; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_28; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_29; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_30; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_31; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_32; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_33; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_34; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_35; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_36; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_37; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_38; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_39; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_40; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_41; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_42; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_43; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_44; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_45; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_46; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_47; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_48; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_49; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_50; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_51; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_52; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_53; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_54; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_55; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_56; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_57; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_58; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_59; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_60; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_61; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_62; // @[CFARCoreWithASR.scala 43:30]
  wire [15:0] laggWindow_io_parallelOut_63; // @[CFARCoreWithASR.scala 43:30]
  wire [6:0] laggWindow_io_cnt; // @[CFARCoreWithASR.scala 43:30]
  wire  laggWindow_io_regFull; // @[CFARCoreWithASR.scala 43:30]
  wire  laggGuard_clock; // @[CFARCoreWithASR.scala 58:29]
  wire  laggGuard_reset; // @[CFARCoreWithASR.scala 58:29]
  wire [3:0] laggGuard_io_depth; // @[CFARCoreWithASR.scala 58:29]
  wire  laggGuard_io_in_ready; // @[CFARCoreWithASR.scala 58:29]
  wire  laggGuard_io_in_valid; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_in_bits; // @[CFARCoreWithASR.scala 58:29]
  wire  laggGuard_io_lastIn; // @[CFARCoreWithASR.scala 58:29]
  wire  laggGuard_io_out_ready; // @[CFARCoreWithASR.scala 58:29]
  wire  laggGuard_io_out_valid; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_out_bits; // @[CFARCoreWithASR.scala 58:29]
  wire  laggGuard_io_lastOut; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_0; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_1; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_2; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_3; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_4; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_5; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_6; // @[CFARCoreWithASR.scala 58:29]
  wire [15:0] laggGuard_io_parallelOut_7; // @[CFARCoreWithASR.scala 58:29]
  wire  cellUnderTest_clock; // @[CFARCoreWithASR.scala 63:29]
  wire  cellUnderTest_reset; // @[CFARCoreWithASR.scala 63:29]
  wire  cellUnderTest_io_in_ready; // @[CFARCoreWithASR.scala 63:29]
  wire  cellUnderTest_io_in_valid; // @[CFARCoreWithASR.scala 63:29]
  wire [15:0] cellUnderTest_io_in_bits; // @[CFARCoreWithASR.scala 63:29]
  wire  cellUnderTest_io_lastIn; // @[CFARCoreWithASR.scala 63:29]
  wire  cellUnderTest_io_out_ready; // @[CFARCoreWithASR.scala 63:29]
  wire  cellUnderTest_io_out_valid; // @[CFARCoreWithASR.scala 63:29]
  wire [15:0] cellUnderTest_io_out_bits; // @[CFARCoreWithASR.scala 63:29]
  wire  cellUnderTest_io_lastOut; // @[CFARCoreWithASR.scala 63:29]
  wire  leadGuard_clock; // @[CFARCoreWithASR.scala 68:25]
  wire  leadGuard_reset; // @[CFARCoreWithASR.scala 68:25]
  wire [3:0] leadGuard_io_depth; // @[CFARCoreWithASR.scala 68:25]
  wire  leadGuard_io_in_ready; // @[CFARCoreWithASR.scala 68:25]
  wire  leadGuard_io_in_valid; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_in_bits; // @[CFARCoreWithASR.scala 68:25]
  wire  leadGuard_io_lastIn; // @[CFARCoreWithASR.scala 68:25]
  wire  leadGuard_io_out_ready; // @[CFARCoreWithASR.scala 68:25]
  wire  leadGuard_io_out_valid; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_out_bits; // @[CFARCoreWithASR.scala 68:25]
  wire  leadGuard_io_lastOut; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_0; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_1; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_2; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_3; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_4; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_5; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_6; // @[CFARCoreWithASR.scala 68:25]
  wire [15:0] leadGuard_io_parallelOut_7; // @[CFARCoreWithASR.scala 68:25]
  wire  leadWindow_clock; // @[CFARCoreWithASR.scala 74:26]
  wire  leadWindow_reset; // @[CFARCoreWithASR.scala 74:26]
  wire [6:0] leadWindow_io_depth; // @[CFARCoreWithASR.scala 74:26]
  wire  leadWindow_io_in_ready; // @[CFARCoreWithASR.scala 74:26]
  wire  leadWindow_io_in_valid; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_in_bits; // @[CFARCoreWithASR.scala 74:26]
  wire  leadWindow_io_lastIn; // @[CFARCoreWithASR.scala 74:26]
  wire  leadWindow_io_out_ready; // @[CFARCoreWithASR.scala 74:26]
  wire  leadWindow_io_out_valid; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_0; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_1; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_2; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_3; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_4; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_5; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_6; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_7; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_8; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_9; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_10; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_11; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_12; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_13; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_14; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_15; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_16; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_17; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_18; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_19; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_20; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_21; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_22; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_23; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_24; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_25; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_26; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_27; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_28; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_29; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_30; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_31; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_32; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_33; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_34; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_35; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_36; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_37; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_38; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_39; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_40; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_41; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_42; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_43; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_44; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_45; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_46; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_47; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_48; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_49; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_50; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_51; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_52; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_53; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_54; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_55; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_56; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_57; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_58; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_59; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_60; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_61; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_62; // @[CFARCoreWithASR.scala 74:26]
  wire [15:0] leadWindow_io_parallelOut_63; // @[CFARCoreWithASR.scala 74:26]
  wire [6:0] leadWindow_io_cnt; // @[CFARCoreWithASR.scala 74:26]
  wire  leadWindow_io_regFull; // @[CFARCoreWithASR.scala 74:26]
  wire  minCircuit_clock; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_0; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_1; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_2; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_3; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_4; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_5; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_6; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_7; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_8; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_9; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_10; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_11; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_12; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_13; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_14; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_in_15; // @[CFARCoreWithASR.scala 207:26]
  wire [4:0] minCircuit_io_inSize; // @[CFARCoreWithASR.scala 207:26]
  wire [19:0] minCircuit_io_out; // @[CFARCoreWithASR.scala 207:26]
  wire  Queue_clock; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_reset; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_io_enq_ready; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_io_enq_valid; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_io_enq_bits_peak; // @[CFARCoreWithASR.scala 417:27]
  wire [15:0] Queue_io_enq_bits_cut; // @[CFARCoreWithASR.scala 417:27]
  wire [15:0] Queue_io_enq_bits_threshold; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_io_deq_ready; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_io_deq_valid; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_io_deq_bits_peak; // @[CFARCoreWithASR.scala 417:27]
  wire [15:0] Queue_io_deq_bits_cut; // @[CFARCoreWithASR.scala 417:27]
  wire [15:0] Queue_io_deq_bits_threshold; // @[CFARCoreWithASR.scala 417:27]
  wire  Queue_1_clock; // @[CFARCoreWithASR.scala 434:27]
  wire  Queue_1_reset; // @[CFARCoreWithASR.scala 434:27]
  wire  Queue_1_io_enq_ready; // @[CFARCoreWithASR.scala 434:27]
  wire  Queue_1_io_enq_valid; // @[CFARCoreWithASR.scala 434:27]
  wire  Queue_1_io_enq_bits; // @[CFARCoreWithASR.scala 434:27]
  wire  Queue_1_io_deq_ready; // @[CFARCoreWithASR.scala 434:27]
  wire  Queue_1_io_deq_valid; // @[CFARCoreWithASR.scala 434:27]
  wire  Queue_1_io_deq_bits; // @[CFARCoreWithASR.scala 434:27]
  wire  _T; // @[CFARCoreWithASR.scala 20:25]
  wire  _T_2; // @[CFARCoreWithASR.scala 20:9]
  wire  _T_3; // @[CFARCoreWithASR.scala 20:9]
  reg  flushing; // @[CFARCoreWithASR.scala 23:25]
  reg [31:0] _RAND_0;
  reg [8:0] cntIn; // @[CFARCoreWithASR.scala 24:22]
  reg [31:0] _RAND_1;
  reg [8:0] cntOut; // @[CFARCoreWithASR.scala 25:23]
  reg [31:0] _RAND_2;
  reg  initialInDone; // @[CFARCoreWithASR.scala 26:30]
  reg [31:0] _RAND_3;
  wire [6:0] _GEN_733; // @[CFARCoreWithASR.scala 37:32]
  wire [7:0] _T_4; // @[CFARCoreWithASR.scala 37:32]
  wire [8:0] latency; // @[CFARCoreWithASR.scala 37:49]
  wire [8:0] _T_5; // @[CFARCoreWithASR.scala 38:26]
  wire [5:0] _T_6; // @[CFARCoreWithASR.scala 38:49]
  wire [8:0] _GEN_734; // @[CFARCoreWithASR.scala 38:43]
  wire [8:0] _T_8; // @[CFARCoreWithASR.scala 38:43]
  wire [8:0] _T_10; // @[CFARCoreWithASR.scala 38:65]
  wire [9:0] _GEN_735; // @[CFARCoreWithASR.scala 38:20]
  wire  _T_11; // @[CFARCoreWithASR.scala 38:20]
  wire  _T_13; // @[CFARCoreWithASR.scala 38:9]
  wire  _T_14; // @[CFARCoreWithASR.scala 38:9]
  reg  lastOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [19:0] sumSubLaggs_0; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_5;
  reg [19:0] sumSubLaggs_1; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_6;
  reg [19:0] sumSubLaggs_2; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_7;
  reg [19:0] sumSubLaggs_3; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_8;
  reg [19:0] sumSubLaggs_4; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_9;
  reg [19:0] sumSubLaggs_5; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_10;
  reg [19:0] sumSubLaggs_6; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_11;
  reg [19:0] sumSubLaggs_7; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_12;
  reg [19:0] sumSubLaggs_8; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_13;
  reg [19:0] sumSubLaggs_9; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_14;
  reg [19:0] sumSubLaggs_10; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_15;
  reg [19:0] sumSubLaggs_11; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_16;
  reg [19:0] sumSubLaggs_12; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_17;
  reg [19:0] sumSubLaggs_13; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_18;
  reg [19:0] sumSubLaggs_14; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_19;
  reg [19:0] sumSubLaggs_15; // @[CFARCoreWithASR.scala 86:28]
  reg [31:0] _RAND_20;
  reg [19:0] sumSubLeads_0; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_21;
  reg [19:0] sumSubLeads_1; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_22;
  reg [19:0] sumSubLeads_2; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_23;
  reg [19:0] sumSubLeads_3; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_24;
  reg [19:0] sumSubLeads_4; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_25;
  reg [19:0] sumSubLeads_5; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_26;
  reg [19:0] sumSubLeads_6; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_27;
  reg [19:0] sumSubLeads_7; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_28;
  reg [19:0] sumSubLeads_8; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_29;
  reg [19:0] sumSubLeads_9; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_30;
  reg [19:0] sumSubLeads_10; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_31;
  reg [19:0] sumSubLeads_11; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_32;
  reg [19:0] sumSubLeads_12; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_33;
  reg [19:0] sumSubLeads_13; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_34;
  reg [19:0] sumSubLeads_14; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_35;
  reg [19:0] sumSubLeads_15; // @[CFARCoreWithASR.scala 87:28]
  reg [31:0] _RAND_36;
  wire  _T_86; // @[CFARCoreWithASR.scala 108:55]
  wire  _T_87; // @[CFARCoreWithASR.scala 108:55]
  wire  _T_88; // @[CFARCoreWithASR.scala 108:55]
  wire  _T_89; // @[CFARCoreWithASR.scala 108:55]
  wire  _T_90; // @[CFARCoreWithASR.scala 108:55]
  wire  _T_92; // @[CFARCoreWithASR.scala 110:58]
  wire  _T_93; // @[CFARCoreWithASR.scala 110:58]
  wire  _T_94; // @[CFARCoreWithASR.scala 110:58]
  wire  _T_95; // @[CFARCoreWithASR.scala 110:58]
  wire  _T_96; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_97; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_98; // @[Mux.scala 87:16]
  wire [15:0] _T_99; // @[Mux.scala 87:16]
  wire [15:0] _T_100; // @[Mux.scala 87:16]
  wire [15:0] _T_101; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg; // @[Mux.scala 87:16]
  wire [15:0] _T_102; // @[Mux.scala 87:16]
  wire [15:0] _T_103; // @[Mux.scala 87:16]
  wire [15:0] _T_104; // @[Mux.scala 87:16]
  wire [15:0] _T_105; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead; // @[Mux.scala 87:16]
  wire [6:0] _T_107; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_108; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_111; // @[CFARCoreWithASR.scala 133:57]
  wire  _T_114; // @[Decoupled.scala 40:37]
  wire  maybeFullLagg_0; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_115; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_736; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_118; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_737; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_121; // @[FixedPointTypeClass.scala 30:68]
  wire  _T_127; // @[Decoupled.scala 40:37]
  wire  _T_128; // @[Decoupled.scala 40:37]
  wire  _T_129; // @[CFARCoreWithASR.scala 170:40]
  wire  maybeFullLead_0; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_130; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_739; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_133; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_740; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_136; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_141; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_145; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_146; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_1; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_1; // @[Mux.scala 87:16]
  wire [6:0] _T_148; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_149; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_152; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_1; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_156; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_742; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_159; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_743; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_162; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_1; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_171; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_745; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_174; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_746; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_177; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_182; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_1; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_188; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_189; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_190; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg_2; // @[Mux.scala 87:16]
  wire [15:0] _T_191; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_2; // @[Mux.scala 87:16]
  wire [6:0] _T_193; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_194; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_197; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_2; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_201; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_748; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_204; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_749; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_207; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_2; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_216; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_751; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_219; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_752; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_222; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_227; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_2; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_231; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_232; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_3; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_3; // @[Mux.scala 87:16]
  wire [6:0] _T_234; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_235; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_238; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_3; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_242; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_754; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_245; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_755; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_248; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_3; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_257; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_757; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_260; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_758; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_263; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_268; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_3; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_276; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_277; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_278; // @[Mux.scala 87:16]
  wire [15:0] _T_279; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg_4; // @[Mux.scala 87:16]
  wire [15:0] _T_280; // @[Mux.scala 87:16]
  wire [15:0] _T_281; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_4; // @[Mux.scala 87:16]
  wire [6:0] _T_283; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_284; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_287; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_4; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_291; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_760; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_294; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_761; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_297; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_4; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_306; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_763; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_309; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_764; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_312; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_317; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_4; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_321; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_322; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_5; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_5; // @[Mux.scala 87:16]
  wire [6:0] _T_324; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_325; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_328; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_5; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_332; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_766; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_335; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_767; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_338; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_5; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_347; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_769; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_350; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_770; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_353; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_358; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_5; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_364; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_365; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_366; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg_6; // @[Mux.scala 87:16]
  wire [15:0] _T_367; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_6; // @[Mux.scala 87:16]
  wire [6:0] _T_369; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_370; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_373; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_6; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_377; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_772; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_380; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_773; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_383; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_6; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_392; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_775; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_395; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_776; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_398; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_403; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_6; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_407; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_408; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_7; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_7; // @[Mux.scala 87:16]
  wire [6:0] _T_410; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_411; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_414; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_7; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_418; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_778; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_421; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_779; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_424; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_7; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_433; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_781; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_436; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_782; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_439; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_444; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_7; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_454; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_455; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_456; // @[Mux.scala 87:16]
  wire [15:0] _T_457; // @[Mux.scala 87:16]
  wire [15:0] _T_458; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg_8; // @[Mux.scala 87:16]
  wire [15:0] _T_459; // @[Mux.scala 87:16]
  wire [15:0] _T_460; // @[Mux.scala 87:16]
  wire [15:0] _T_461; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_8; // @[Mux.scala 87:16]
  wire [6:0] _T_463; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_464; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_467; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_8; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_471; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_784; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_474; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_785; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_477; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_8; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_486; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_787; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_489; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_788; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_492; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_497; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_8; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_501; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_502; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_9; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_9; // @[Mux.scala 87:16]
  wire [6:0] _T_504; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_505; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_508; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_9; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_512; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_790; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_515; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_791; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_518; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_9; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_527; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_793; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_530; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_794; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_533; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_538; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_9; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_544; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_545; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_546; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg_10; // @[Mux.scala 87:16]
  wire [15:0] _T_547; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_10; // @[Mux.scala 87:16]
  wire [6:0] _T_549; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_550; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_553; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_10; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_557; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_796; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_560; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_797; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_563; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_10; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_572; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_799; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_575; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_800; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_578; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_583; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_10; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_587; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_588; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_11; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_11; // @[Mux.scala 87:16]
  wire [6:0] _T_590; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_591; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_594; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_11; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_598; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_802; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_601; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_803; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_604; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_11; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_613; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_805; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_616; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_806; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_619; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_624; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_11; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_632; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_633; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_634; // @[Mux.scala 87:16]
  wire [15:0] _T_635; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg_12; // @[Mux.scala 87:16]
  wire [15:0] _T_636; // @[Mux.scala 87:16]
  wire [15:0] _T_637; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_12; // @[Mux.scala 87:16]
  wire [6:0] _T_639; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_640; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_643; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_12; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_647; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_808; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_650; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_809; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_653; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_12; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_662; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_811; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_665; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_812; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_668; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_673; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_12; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_677; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_678; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_13; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_13; // @[Mux.scala 87:16]
  wire [6:0] _T_680; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_681; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_684; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_13; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_688; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_814; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_691; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_815; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_694; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_13; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_703; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_817; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_706; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_818; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_709; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_714; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_13; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_720; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_721; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] _T_722; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLagg_14; // @[Mux.scala 87:16]
  wire [15:0] _T_723; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_14; // @[Mux.scala 87:16]
  wire [6:0] _T_725; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_726; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_729; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_14; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_733; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_820; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_736; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_821; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_739; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_14; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_748; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_823; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_751; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_824; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_754; // @[FixedPointTypeClass.scala 30:68]
  wire [6:0] _T_759; // @[CFARCoreWithASR.scala 103:76]
  wire [6:0] endIndex_14; // @[CFARCoreWithASR.scala 103:94]
  wire  _T_763; // @[CFARCoreWithASR.scala 110:76]
  wire  _T_764; // @[CFARCoreWithASR.scala 110:64]
  wire [15:0] minusOperandLagg_15; // @[Mux.scala 87:16]
  wire [15:0] minusOperandLead_15; // @[Mux.scala 87:16]
  wire [6:0] _T_766; // @[CFARCoreWithASR.scala 132:69]
  wire  _T_767; // @[CFARCoreWithASR.scala 132:57]
  wire  _T_770; // @[CFARCoreWithASR.scala 133:57]
  wire  maybeFullLagg_15; // @[CFARCoreWithASR.scala 133:32]
  wire  _T_774; // @[CFARCoreWithASR.scala 147:35]
  wire [19:0] _GEN_826; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_777; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_827; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_780; // @[FixedPointTypeClass.scala 30:68]
  wire  maybeFullLead_15; // @[CFARCoreWithASR.scala 132:32]
  wire  _T_789; // @[CFARCoreWithASR.scala 172:35]
  wire [19:0] _GEN_829; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_792; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _GEN_830; // @[FixedPointTypeClass.scala 30:68]
  wire [19:0] _T_795; // @[FixedPointTypeClass.scala 30:68]
  wire  _T_801; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_804; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_808; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_809; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_810; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_811; // @[Cat.scala 29:58]
  wire [2:0] diffInSubSize; // @[CFARCoreWithASR.scala 193:45]
  wire  _T_814; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_0; // @[Order.scala 56:31]
  wire  _T_815; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_1; // @[Order.scala 56:31]
  wire  _T_816; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_2; // @[Order.scala 56:31]
  wire  _T_817; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_3; // @[Order.scala 56:31]
  wire  _T_818; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_4; // @[Order.scala 56:31]
  wire  _T_819; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_5; // @[Order.scala 56:31]
  wire  _T_820; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_6; // @[Order.scala 56:31]
  wire  _T_821; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_7; // @[Order.scala 56:31]
  wire  _T_822; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_8; // @[Order.scala 56:31]
  wire  _T_823; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_9; // @[Order.scala 56:31]
  wire  _T_824; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_10; // @[Order.scala 56:31]
  wire  _T_825; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_11; // @[Order.scala 56:31]
  wire  _T_826; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_12; // @[Order.scala 56:31]
  wire  _T_827; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_13; // @[Order.scala 56:31]
  wire  _T_828; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_14; // @[Order.scala 56:31]
  wire  _T_829; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] max_15; // @[Order.scala 56:31]
  wire  activeSums_0; // @[CFARCoreWithASR.scala 110:29]
  wire  _T_864; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_127; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_128; // @[CFARCoreWithASR.scala 202:27]
  wire [1:0] _GEN_832; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_129; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_130; // @[CFARCoreWithASR.scala 202:27]
  wire [2:0] _GEN_834; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_131; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_132; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_133; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_134; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_838; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_135; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_136; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_137; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_138; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_139; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_140; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_141; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_142; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_143; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_144; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_145; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_146; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_147; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_148; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_149; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_150; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_151; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_152; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_153; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_154; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_155; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_156; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_157; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_158; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_1; // @[CFARCoreWithASR.scala 110:29]
  wire  _T_866; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_159; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_160; // @[CFARCoreWithASR.scala 202:27]
  wire [1:0] _GEN_846; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_161; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_162; // @[CFARCoreWithASR.scala 202:27]
  wire [2:0] _GEN_848; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_163; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_164; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_165; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_166; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_852; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_167; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_168; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_169; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_170; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_171; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_172; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_173; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_174; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_175; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_176; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_177; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_178; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_179; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_180; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_181; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_182; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_183; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_184; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_185; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_186; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_187; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_188; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_189; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_190; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_2; // @[CFARCoreWithASR.scala 110:29]
  wire [1:0] _T_868; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_191; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_192; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_193; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_194; // @[CFARCoreWithASR.scala 202:27]
  wire [2:0] _GEN_860; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_195; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_196; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_197; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_198; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_864; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_199; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_200; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_201; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_202; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_203; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_204; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_205; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_206; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_207; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_208; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_209; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_210; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_211; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_212; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_213; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_214; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_215; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_216; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_217; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_218; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_219; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_220; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_221; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_222; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_3; // @[CFARCoreWithASR.scala 110:29]
  wire [1:0] _T_870; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_223; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_224; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_225; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_226; // @[CFARCoreWithASR.scala 202:27]
  wire [2:0] _GEN_872; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_227; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_228; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_229; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_230; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_876; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_231; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_232; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_233; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_234; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_235; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_236; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_237; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_238; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_239; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_240; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_241; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_242; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_243; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_244; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_245; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_246; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_247; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_248; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_249; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_250; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_251; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_252; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_253; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_254; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_4; // @[CFARCoreWithASR.scala 110:29]
  wire [2:0] _T_872; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_255; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_256; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_257; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_258; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_259; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_260; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_261; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_262; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_884; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_263; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_264; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_265; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_266; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_267; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_268; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_269; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_270; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_271; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_272; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_273; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_274; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_275; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_276; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_277; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_278; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_279; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_280; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_281; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_282; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_283; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_284; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_285; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_286; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_5; // @[CFARCoreWithASR.scala 110:29]
  wire [2:0] _T_874; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_287; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_288; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_289; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_290; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_291; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_292; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_293; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_294; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_892; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_295; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_296; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_297; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_298; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_299; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_300; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_301; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_302; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_303; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_304; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_305; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_306; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_307; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_308; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_309; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_310; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_311; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_312; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_313; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_314; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_315; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_316; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_317; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_318; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_6; // @[CFARCoreWithASR.scala 110:29]
  wire [2:0] _T_876; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_319; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_320; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_321; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_322; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_323; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_324; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_325; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_326; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_900; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_327; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_328; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_329; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_330; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_331; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_332; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_333; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_334; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_335; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_336; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_337; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_338; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_339; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_340; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_341; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_342; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_343; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_344; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_345; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_346; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_347; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_348; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_349; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_350; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_7; // @[CFARCoreWithASR.scala 110:29]
  wire [2:0] _T_878; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_351; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_352; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_353; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_354; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_355; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_356; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_357; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_358; // @[CFARCoreWithASR.scala 202:27]
  wire [3:0] _GEN_908; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_359; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_360; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_361; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_362; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_363; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_364; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_365; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_366; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_367; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_368; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_369; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_370; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_371; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_372; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_373; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_374; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_375; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_376; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_377; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_378; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_379; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_380; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_381; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_382; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_8; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_880; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_383; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_384; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_385; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_386; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_387; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_388; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_389; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_390; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_391; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_392; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_393; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_394; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_395; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_396; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_397; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_398; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_399; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_400; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_401; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_402; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_403; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_404; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_405; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_406; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_407; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_408; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_409; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_410; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_411; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_412; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_413; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_414; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_9; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_882; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_415; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_416; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_417; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_418; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_419; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_420; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_421; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_422; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_423; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_424; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_425; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_426; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_427; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_428; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_429; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_430; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_431; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_432; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_433; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_434; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_435; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_436; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_437; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_438; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_439; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_440; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_441; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_442; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_443; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_444; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_445; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_446; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_10; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_884; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_447; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_448; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_449; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_450; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_451; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_452; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_453; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_454; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_455; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_456; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_457; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_458; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_459; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_460; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_461; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_462; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_463; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_464; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_465; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_466; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_467; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_468; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_469; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_470; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_471; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_472; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_473; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_474; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_475; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_476; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_477; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_478; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_11; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_886; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_479; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_480; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_481; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_482; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_483; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_484; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_485; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_486; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_487; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_488; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_489; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_490; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_491; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_492; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_493; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_494; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_495; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_496; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_497; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_498; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_499; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_500; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_501; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_502; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_503; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_504; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_505; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_506; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_507; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_508; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_509; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_510; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_12; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_888; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_511; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_512; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_513; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_514; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_515; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_516; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_517; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_518; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_519; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_520; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_521; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_522; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_523; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_524; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_525; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_526; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_527; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_528; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_529; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_530; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_531; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_532; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_533; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_534; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_535; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_536; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_537; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_538; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_539; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_540; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_541; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_542; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_13; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_890; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_543; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_544; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_545; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_546; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_547; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_548; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_549; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_550; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_551; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_552; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_553; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_554; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_555; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_556; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_557; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_558; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_559; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_560; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_561; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_562; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_563; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_564; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_565; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_566; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_567; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_568; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_569; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_570; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_571; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_572; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_573; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_574; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_14; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_892; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_575; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_576; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_577; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_578; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_579; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_580; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_581; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_582; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_583; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_584; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_585; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_586; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_587; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_588; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_589; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_590; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_591; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_592; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_593; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_594; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_595; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_596; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_597; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_598; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_599; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_600; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_601; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_602; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_603; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_604; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_605; // @[CFARCoreWithASR.scala 200:32]
  wire [19:0] _GEN_606; // @[CFARCoreWithASR.scala 200:32]
  wire  activeSums_15; // @[CFARCoreWithASR.scala 110:29]
  wire [3:0] _T_894; // @[CFARCoreWithASR.scala 201:29]
  wire [19:0] _GEN_607; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_608; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_609; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_610; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_611; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_612; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_613; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_614; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_615; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_616; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_617; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_618; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_619; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_620; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_621; // @[CFARCoreWithASR.scala 202:27]
  wire [19:0] _GEN_622; // @[CFARCoreWithASR.scala 202:27]
  wire [6:0] _T_908; // @[CFARCoreWithASR.scala 209:46]
  wire [19:0] clutterRepr; // @[FixedPointTypeClass.scala 118:51]
  wire [8:0] _T_924; // @[CFARCoreWithASR.scala 216:20]
  wire [8:0] _T_926; // @[CFARCoreWithASR.scala 218:28]
  wire  _T_927; // @[CFARCoreWithASR.scala 218:15]
  wire  _T_929; // @[CFARCoreWithASR.scala 218:35]
  wire  _GEN_640; // @[CFARCoreWithASR.scala 218:52]
  wire  _T_930; // @[Decoupled.scala 40:37]
  wire  _T_931; // @[CFARCoreWithASR.scala 222:20]
  wire [8:0] _T_934; // @[CFARCoreWithASR.scala 226:22]
  wire [9:0] _T_936; // @[CFARCoreWithASR.scala 228:31]
  wire [9:0] _GEN_916; // @[CFARCoreWithASR.scala 228:16]
  wire  _T_937; // @[CFARCoreWithASR.scala 228:16]
  wire  _T_939; // @[CFARCoreWithASR.scala 228:38]
  wire  _T_942; // @[CFARCoreWithASR.scala 228:55]
  wire  _GEN_644; // @[CFARCoreWithASR.scala 232:20]
  reg  flushingDelayed; // @[CFARUtils.scala 286:20]
  reg [31:0] _RAND_37;
  wire [19:0] leftThr; // @[FixedPointTypeClass.scala 118:51]
  wire [19:0] rightThr; // @[FixedPointTypeClass.scala 118:51]
  wire  _T_944; // @[FixedPointTypeClass.scala 55:59]
  wire [19:0] greatestOf; // @[CFARCoreWithASR.scala 289:23]
  wire  _T_945; // @[FixedPointTypeClass.scala 53:59]
  wire [19:0] smallestOf; // @[CFARCoreWithASR.scala 290:23]
  wire [19:0] _T_948; // @[FixedPointTypeClass.scala 20:58]
  wire [18:0] _T_949; // @[FixedPointTypeClass.scala 117:50]
  wire  _T_950; // @[Mux.scala 68:19]
  wire [19:0] _T_951; // @[Mux.scala 68:16]
  wire  _T_952; // @[Mux.scala 68:19]
  wire [19:0] _T_953; // @[Mux.scala 68:16]
  wire  _T_954; // @[Mux.scala 68:19]
  wire [19:0] _T_955; // @[Mux.scala 68:16]
  wire  _T_956; // @[Mux.scala 68:19]
  wire [19:0] thrByModes; // @[Mux.scala 68:16]
  reg  enableRightThr; // @[CFARCoreWithASR.scala 299:31]
  reg [31:0] _RAND_38;
  wire  _T_957; // @[CFARCoreWithASR.scala 300:9]
  wire  _T_958; // @[Decoupled.scala 40:37]
  wire  _T_959; // @[CFARCoreWithASR.scala 300:34]
  wire  _GEN_651; // @[CFARCoreWithASR.scala 300:63]
  wire  _T_960; // @[CFARCoreWithASR.scala 313:50]
  wire  _T_961; // @[CFARCoreWithASR.scala 315:60]
  wire  _T_962; // @[CFARCoreWithASR.scala 315:57]
  wire [19:0] _T_963; // @[CFARCoreWithASR.scala 315:87]
  wire [19:0] _T_964; // @[CFARCoreWithASR.scala 315:41]
  wire [19:0] thrWithoutScaling; // @[CFARCoreWithASR.scala 313:27]
  wire [19:0] _GEN_917; // @[FixedPointTypeClass.scala 211:35]
  reg [35:0] _T_966; // @[Reg.scala 15:16]
  reg [63:0] _RAND_39;
  wire [22:0] threshold; // @[FixedPointTypeClass.scala 153:43]
  reg [15:0] cutDelayed; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  wire  _T_967; // @[CFARCoreWithASR.scala 394:53]
  wire [6:0] _T_969; // @[CFARCoreWithASR.scala 394:103]
  wire [3:0] _T_972; // @[CFARCoreWithASR.scala 394:150]
  wire [15:0] _GEN_655; // @[CFARCoreWithASR.scala 394:38]
  wire [15:0] _GEN_719; // @[CFARCoreWithASR.scala 394:38]
  reg [15:0] leftNeighb; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [15:0] rightNeighb; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  wire  _T_977; // @[FixedPointTypeClass.scala 55:59]
  wire  _T_978; // @[FixedPointTypeClass.scala 55:59]
  wire  isLocalMax; // @[CFARCoreWithASR.scala 396:44]
  wire [16:0] _GEN_918; // @[FixedPointTypeClass.scala 55:59]
  wire [22:0] _GEN_919; // @[FixedPointTypeClass.scala 55:59]
  wire  isPeak; // @[FixedPointTypeClass.scala 55:59]
  wire  _T_979; // @[CFARCoreWithASR.scala 418:20]
  wire  _T_980; // @[CFARCoreWithASR.scala 418:54]
  wire  _T_981; // @[CFARCoreWithASR.scala 418:51]
  reg  _T_985; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg  _T_986; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  wire  _T_987; // @[CFARCoreWithASR.scala 419:121]
  wire  _T_989; // @[CFARCoreWithASR.scala 430:65]
  reg  _T_993; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg  _T_994; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  wire  _T_995; // @[CFARCoreWithASR.scala 435:121]
  wire [21:0] _GEN_921; // @[CFARCoreWithASR.scala 423:37]
  AdjustableShiftRegisterStream laggWindow ( // @[CFARCoreWithASR.scala 43:30]
    .clock(laggWindow_clock),
    .reset(laggWindow_reset),
    .io_depth(laggWindow_io_depth),
    .io_in_ready(laggWindow_io_in_ready),
    .io_in_valid(laggWindow_io_in_valid),
    .io_in_bits(laggWindow_io_in_bits),
    .io_lastIn(laggWindow_io_lastIn),
    .io_out_ready(laggWindow_io_out_ready),
    .io_out_valid(laggWindow_io_out_valid),
    .io_out_bits(laggWindow_io_out_bits),
    .io_lastOut(laggWindow_io_lastOut),
    .io_parallelOut_0(laggWindow_io_parallelOut_0),
    .io_parallelOut_1(laggWindow_io_parallelOut_1),
    .io_parallelOut_2(laggWindow_io_parallelOut_2),
    .io_parallelOut_3(laggWindow_io_parallelOut_3),
    .io_parallelOut_4(laggWindow_io_parallelOut_4),
    .io_parallelOut_5(laggWindow_io_parallelOut_5),
    .io_parallelOut_6(laggWindow_io_parallelOut_6),
    .io_parallelOut_7(laggWindow_io_parallelOut_7),
    .io_parallelOut_8(laggWindow_io_parallelOut_8),
    .io_parallelOut_9(laggWindow_io_parallelOut_9),
    .io_parallelOut_10(laggWindow_io_parallelOut_10),
    .io_parallelOut_11(laggWindow_io_parallelOut_11),
    .io_parallelOut_12(laggWindow_io_parallelOut_12),
    .io_parallelOut_13(laggWindow_io_parallelOut_13),
    .io_parallelOut_14(laggWindow_io_parallelOut_14),
    .io_parallelOut_15(laggWindow_io_parallelOut_15),
    .io_parallelOut_16(laggWindow_io_parallelOut_16),
    .io_parallelOut_17(laggWindow_io_parallelOut_17),
    .io_parallelOut_18(laggWindow_io_parallelOut_18),
    .io_parallelOut_19(laggWindow_io_parallelOut_19),
    .io_parallelOut_20(laggWindow_io_parallelOut_20),
    .io_parallelOut_21(laggWindow_io_parallelOut_21),
    .io_parallelOut_22(laggWindow_io_parallelOut_22),
    .io_parallelOut_23(laggWindow_io_parallelOut_23),
    .io_parallelOut_24(laggWindow_io_parallelOut_24),
    .io_parallelOut_25(laggWindow_io_parallelOut_25),
    .io_parallelOut_26(laggWindow_io_parallelOut_26),
    .io_parallelOut_27(laggWindow_io_parallelOut_27),
    .io_parallelOut_28(laggWindow_io_parallelOut_28),
    .io_parallelOut_29(laggWindow_io_parallelOut_29),
    .io_parallelOut_30(laggWindow_io_parallelOut_30),
    .io_parallelOut_31(laggWindow_io_parallelOut_31),
    .io_parallelOut_32(laggWindow_io_parallelOut_32),
    .io_parallelOut_33(laggWindow_io_parallelOut_33),
    .io_parallelOut_34(laggWindow_io_parallelOut_34),
    .io_parallelOut_35(laggWindow_io_parallelOut_35),
    .io_parallelOut_36(laggWindow_io_parallelOut_36),
    .io_parallelOut_37(laggWindow_io_parallelOut_37),
    .io_parallelOut_38(laggWindow_io_parallelOut_38),
    .io_parallelOut_39(laggWindow_io_parallelOut_39),
    .io_parallelOut_40(laggWindow_io_parallelOut_40),
    .io_parallelOut_41(laggWindow_io_parallelOut_41),
    .io_parallelOut_42(laggWindow_io_parallelOut_42),
    .io_parallelOut_43(laggWindow_io_parallelOut_43),
    .io_parallelOut_44(laggWindow_io_parallelOut_44),
    .io_parallelOut_45(laggWindow_io_parallelOut_45),
    .io_parallelOut_46(laggWindow_io_parallelOut_46),
    .io_parallelOut_47(laggWindow_io_parallelOut_47),
    .io_parallelOut_48(laggWindow_io_parallelOut_48),
    .io_parallelOut_49(laggWindow_io_parallelOut_49),
    .io_parallelOut_50(laggWindow_io_parallelOut_50),
    .io_parallelOut_51(laggWindow_io_parallelOut_51),
    .io_parallelOut_52(laggWindow_io_parallelOut_52),
    .io_parallelOut_53(laggWindow_io_parallelOut_53),
    .io_parallelOut_54(laggWindow_io_parallelOut_54),
    .io_parallelOut_55(laggWindow_io_parallelOut_55),
    .io_parallelOut_56(laggWindow_io_parallelOut_56),
    .io_parallelOut_57(laggWindow_io_parallelOut_57),
    .io_parallelOut_58(laggWindow_io_parallelOut_58),
    .io_parallelOut_59(laggWindow_io_parallelOut_59),
    .io_parallelOut_60(laggWindow_io_parallelOut_60),
    .io_parallelOut_61(laggWindow_io_parallelOut_61),
    .io_parallelOut_62(laggWindow_io_parallelOut_62),
    .io_parallelOut_63(laggWindow_io_parallelOut_63),
    .io_cnt(laggWindow_io_cnt),
    .io_regFull(laggWindow_io_regFull)
  );
  AdjustableShiftRegisterStream_1 laggGuard ( // @[CFARCoreWithASR.scala 58:29]
    .clock(laggGuard_clock),
    .reset(laggGuard_reset),
    .io_depth(laggGuard_io_depth),
    .io_in_ready(laggGuard_io_in_ready),
    .io_in_valid(laggGuard_io_in_valid),
    .io_in_bits(laggGuard_io_in_bits),
    .io_lastIn(laggGuard_io_lastIn),
    .io_out_ready(laggGuard_io_out_ready),
    .io_out_valid(laggGuard_io_out_valid),
    .io_out_bits(laggGuard_io_out_bits),
    .io_lastOut(laggGuard_io_lastOut),
    .io_parallelOut_0(laggGuard_io_parallelOut_0),
    .io_parallelOut_1(laggGuard_io_parallelOut_1),
    .io_parallelOut_2(laggGuard_io_parallelOut_2),
    .io_parallelOut_3(laggGuard_io_parallelOut_3),
    .io_parallelOut_4(laggGuard_io_parallelOut_4),
    .io_parallelOut_5(laggGuard_io_parallelOut_5),
    .io_parallelOut_6(laggGuard_io_parallelOut_6),
    .io_parallelOut_7(laggGuard_io_parallelOut_7)
  );
  CellUnderTest cellUnderTest ( // @[CFARCoreWithASR.scala 63:29]
    .clock(cellUnderTest_clock),
    .reset(cellUnderTest_reset),
    .io_in_ready(cellUnderTest_io_in_ready),
    .io_in_valid(cellUnderTest_io_in_valid),
    .io_in_bits(cellUnderTest_io_in_bits),
    .io_lastIn(cellUnderTest_io_lastIn),
    .io_out_ready(cellUnderTest_io_out_ready),
    .io_out_valid(cellUnderTest_io_out_valid),
    .io_out_bits(cellUnderTest_io_out_bits),
    .io_lastOut(cellUnderTest_io_lastOut)
  );
  AdjustableShiftRegisterStream_1 leadGuard ( // @[CFARCoreWithASR.scala 68:25]
    .clock(leadGuard_clock),
    .reset(leadGuard_reset),
    .io_depth(leadGuard_io_depth),
    .io_in_ready(leadGuard_io_in_ready),
    .io_in_valid(leadGuard_io_in_valid),
    .io_in_bits(leadGuard_io_in_bits),
    .io_lastIn(leadGuard_io_lastIn),
    .io_out_ready(leadGuard_io_out_ready),
    .io_out_valid(leadGuard_io_out_valid),
    .io_out_bits(leadGuard_io_out_bits),
    .io_lastOut(leadGuard_io_lastOut),
    .io_parallelOut_0(leadGuard_io_parallelOut_0),
    .io_parallelOut_1(leadGuard_io_parallelOut_1),
    .io_parallelOut_2(leadGuard_io_parallelOut_2),
    .io_parallelOut_3(leadGuard_io_parallelOut_3),
    .io_parallelOut_4(leadGuard_io_parallelOut_4),
    .io_parallelOut_5(leadGuard_io_parallelOut_5),
    .io_parallelOut_6(leadGuard_io_parallelOut_6),
    .io_parallelOut_7(leadGuard_io_parallelOut_7)
  );
  AdjustableShiftRegisterStream_3 leadWindow ( // @[CFARCoreWithASR.scala 74:26]
    .clock(leadWindow_clock),
    .reset(leadWindow_reset),
    .io_depth(leadWindow_io_depth),
    .io_in_ready(leadWindow_io_in_ready),
    .io_in_valid(leadWindow_io_in_valid),
    .io_in_bits(leadWindow_io_in_bits),
    .io_lastIn(leadWindow_io_lastIn),
    .io_out_ready(leadWindow_io_out_ready),
    .io_out_valid(leadWindow_io_out_valid),
    .io_parallelOut_0(leadWindow_io_parallelOut_0),
    .io_parallelOut_1(leadWindow_io_parallelOut_1),
    .io_parallelOut_2(leadWindow_io_parallelOut_2),
    .io_parallelOut_3(leadWindow_io_parallelOut_3),
    .io_parallelOut_4(leadWindow_io_parallelOut_4),
    .io_parallelOut_5(leadWindow_io_parallelOut_5),
    .io_parallelOut_6(leadWindow_io_parallelOut_6),
    .io_parallelOut_7(leadWindow_io_parallelOut_7),
    .io_parallelOut_8(leadWindow_io_parallelOut_8),
    .io_parallelOut_9(leadWindow_io_parallelOut_9),
    .io_parallelOut_10(leadWindow_io_parallelOut_10),
    .io_parallelOut_11(leadWindow_io_parallelOut_11),
    .io_parallelOut_12(leadWindow_io_parallelOut_12),
    .io_parallelOut_13(leadWindow_io_parallelOut_13),
    .io_parallelOut_14(leadWindow_io_parallelOut_14),
    .io_parallelOut_15(leadWindow_io_parallelOut_15),
    .io_parallelOut_16(leadWindow_io_parallelOut_16),
    .io_parallelOut_17(leadWindow_io_parallelOut_17),
    .io_parallelOut_18(leadWindow_io_parallelOut_18),
    .io_parallelOut_19(leadWindow_io_parallelOut_19),
    .io_parallelOut_20(leadWindow_io_parallelOut_20),
    .io_parallelOut_21(leadWindow_io_parallelOut_21),
    .io_parallelOut_22(leadWindow_io_parallelOut_22),
    .io_parallelOut_23(leadWindow_io_parallelOut_23),
    .io_parallelOut_24(leadWindow_io_parallelOut_24),
    .io_parallelOut_25(leadWindow_io_parallelOut_25),
    .io_parallelOut_26(leadWindow_io_parallelOut_26),
    .io_parallelOut_27(leadWindow_io_parallelOut_27),
    .io_parallelOut_28(leadWindow_io_parallelOut_28),
    .io_parallelOut_29(leadWindow_io_parallelOut_29),
    .io_parallelOut_30(leadWindow_io_parallelOut_30),
    .io_parallelOut_31(leadWindow_io_parallelOut_31),
    .io_parallelOut_32(leadWindow_io_parallelOut_32),
    .io_parallelOut_33(leadWindow_io_parallelOut_33),
    .io_parallelOut_34(leadWindow_io_parallelOut_34),
    .io_parallelOut_35(leadWindow_io_parallelOut_35),
    .io_parallelOut_36(leadWindow_io_parallelOut_36),
    .io_parallelOut_37(leadWindow_io_parallelOut_37),
    .io_parallelOut_38(leadWindow_io_parallelOut_38),
    .io_parallelOut_39(leadWindow_io_parallelOut_39),
    .io_parallelOut_40(leadWindow_io_parallelOut_40),
    .io_parallelOut_41(leadWindow_io_parallelOut_41),
    .io_parallelOut_42(leadWindow_io_parallelOut_42),
    .io_parallelOut_43(leadWindow_io_parallelOut_43),
    .io_parallelOut_44(leadWindow_io_parallelOut_44),
    .io_parallelOut_45(leadWindow_io_parallelOut_45),
    .io_parallelOut_46(leadWindow_io_parallelOut_46),
    .io_parallelOut_47(leadWindow_io_parallelOut_47),
    .io_parallelOut_48(leadWindow_io_parallelOut_48),
    .io_parallelOut_49(leadWindow_io_parallelOut_49),
    .io_parallelOut_50(leadWindow_io_parallelOut_50),
    .io_parallelOut_51(leadWindow_io_parallelOut_51),
    .io_parallelOut_52(leadWindow_io_parallelOut_52),
    .io_parallelOut_53(leadWindow_io_parallelOut_53),
    .io_parallelOut_54(leadWindow_io_parallelOut_54),
    .io_parallelOut_55(leadWindow_io_parallelOut_55),
    .io_parallelOut_56(leadWindow_io_parallelOut_56),
    .io_parallelOut_57(leadWindow_io_parallelOut_57),
    .io_parallelOut_58(leadWindow_io_parallelOut_58),
    .io_parallelOut_59(leadWindow_io_parallelOut_59),
    .io_parallelOut_60(leadWindow_io_parallelOut_60),
    .io_parallelOut_61(leadWindow_io_parallelOut_61),
    .io_parallelOut_62(leadWindow_io_parallelOut_62),
    .io_parallelOut_63(leadWindow_io_parallelOut_63),
    .io_cnt(leadWindow_io_cnt),
    .io_regFull(leadWindow_io_regFull)
  );
  MinimumCircuit minCircuit ( // @[CFARCoreWithASR.scala 207:26]
    .clock(minCircuit_clock),
    .io_in_0(minCircuit_io_in_0),
    .io_in_1(minCircuit_io_in_1),
    .io_in_2(minCircuit_io_in_2),
    .io_in_3(minCircuit_io_in_3),
    .io_in_4(minCircuit_io_in_4),
    .io_in_5(minCircuit_io_in_5),
    .io_in_6(minCircuit_io_in_6),
    .io_in_7(minCircuit_io_in_7),
    .io_in_8(minCircuit_io_in_8),
    .io_in_9(minCircuit_io_in_9),
    .io_in_10(minCircuit_io_in_10),
    .io_in_11(minCircuit_io_in_11),
    .io_in_12(minCircuit_io_in_12),
    .io_in_13(minCircuit_io_in_13),
    .io_in_14(minCircuit_io_in_14),
    .io_in_15(minCircuit_io_in_15),
    .io_inSize(minCircuit_io_inSize),
    .io_out(minCircuit_io_out)
  );
  Queue_5 Queue ( // @[CFARCoreWithASR.scala 417:27]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_peak(Queue_io_enq_bits_peak),
    .io_enq_bits_cut(Queue_io_enq_bits_cut),
    .io_enq_bits_threshold(Queue_io_enq_bits_threshold),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_peak(Queue_io_deq_bits_peak),
    .io_deq_bits_cut(Queue_io_deq_bits_cut),
    .io_deq_bits_threshold(Queue_io_deq_bits_threshold)
  );
  Queue_6 Queue_1 ( // @[CFARCoreWithASR.scala 434:27]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  assign _T = io_windowCells >= io_subCells; // @[CFARCoreWithASR.scala 20:25]
  assign _T_2 = _T | reset; // @[CFARCoreWithASR.scala 20:9]
  assign _T_3 = ~_T_2; // @[CFARCoreWithASR.scala 20:9]
  assign _GEN_733 = {{3'd0}, io_guardCells}; // @[CFARCoreWithASR.scala 37:32]
  assign _T_4 = io_windowCells + _GEN_733; // @[CFARCoreWithASR.scala 37:32]
  assign latency = _T_4 + 8'h1; // @[CFARCoreWithASR.scala 37:49]
  assign _T_5 = 7'h2 * io_windowCells; // @[CFARCoreWithASR.scala 38:26]
  assign _T_6 = 4'h2 * io_guardCells; // @[CFARCoreWithASR.scala 38:49]
  assign _GEN_734 = {{3'd0}, _T_6}; // @[CFARCoreWithASR.scala 38:43]
  assign _T_8 = _T_5 + _GEN_734; // @[CFARCoreWithASR.scala 38:43]
  assign _T_10 = _T_8 + 9'h1; // @[CFARCoreWithASR.scala 38:65]
  assign _GEN_735 = {{1'd0}, _T_10}; // @[CFARCoreWithASR.scala 38:20]
  assign _T_11 = io_fftWin > _GEN_735; // @[CFARCoreWithASR.scala 38:20]
  assign _T_13 = _T_11 | reset; // @[CFARCoreWithASR.scala 38:9]
  assign _T_14 = ~_T_13; // @[CFARCoreWithASR.scala 38:9]
  assign _T_86 = 7'h4 == io_subCells; // @[CFARCoreWithASR.scala 108:55]
  assign _T_87 = 7'h8 == io_subCells; // @[CFARCoreWithASR.scala 108:55]
  assign _T_88 = 7'h10 == io_subCells; // @[CFARCoreWithASR.scala 108:55]
  assign _T_89 = 7'h20 == io_subCells; // @[CFARCoreWithASR.scala 108:55]
  assign _T_90 = 7'h40 == io_subCells; // @[CFARCoreWithASR.scala 108:55]
  assign _T_92 = _T_86 | _T_87; // @[CFARCoreWithASR.scala 110:58]
  assign _T_93 = _T_92 | _T_88; // @[CFARCoreWithASR.scala 110:58]
  assign _T_94 = _T_93 | _T_89; // @[CFARCoreWithASR.scala 110:58]
  assign _T_95 = _T_94 | _T_90; // @[CFARCoreWithASR.scala 110:58]
  assign _T_96 = io_subCells <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_97 = _T_95 & _T_96; // @[CFARCoreWithASR.scala 110:64]
  assign _T_98 = _T_90 ? $signed(laggWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_99 = _T_89 ? $signed(laggWindow_io_parallelOut_31) : $signed(_T_98); // @[Mux.scala 87:16]
  assign _T_100 = _T_88 ? $signed(laggWindow_io_parallelOut_15) : $signed(_T_99); // @[Mux.scala 87:16]
  assign _T_101 = _T_87 ? $signed(laggWindow_io_parallelOut_7) : $signed(_T_100); // @[Mux.scala 87:16]
  assign minusOperandLagg = _T_86 ? $signed(laggWindow_io_parallelOut_3) : $signed(_T_101); // @[Mux.scala 87:16]
  assign _T_102 = _T_90 ? $signed(leadWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_103 = _T_89 ? $signed(leadWindow_io_parallelOut_31) : $signed(_T_102); // @[Mux.scala 87:16]
  assign _T_104 = _T_88 ? $signed(leadWindow_io_parallelOut_15) : $signed(_T_103); // @[Mux.scala 87:16]
  assign _T_105 = _T_87 ? $signed(leadWindow_io_parallelOut_7) : $signed(_T_104); // @[Mux.scala 87:16]
  assign minusOperandLead = _T_86 ? $signed(leadWindow_io_parallelOut_3) : $signed(_T_105); // @[Mux.scala 87:16]
  assign _T_107 = io_subCells - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_108 = leadWindow_io_cnt > _T_107; // @[CFARCoreWithASR.scala 132:57]
  assign _T_111 = laggWindow_io_cnt > _T_107; // @[CFARCoreWithASR.scala 133:57]
  assign _T_114 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign maybeFullLagg_0 = _T_111; // @[CFARCoreWithASR.scala 133:32]
  assign _T_115 = laggWindow_io_regFull | maybeFullLagg_0; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_736 = {{4{laggWindow_io_in_bits[15]}},laggWindow_io_in_bits}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_118 = $signed(sumSubLaggs_0) + $signed(_GEN_736); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_737 = {{4{minusOperandLagg[15]}},minusOperandLagg}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_121 = $signed(_T_118) - $signed(_GEN_737); // @[FixedPointTypeClass.scala 30:68]
  assign _T_127 = leadWindow_io_in_ready & leadWindow_io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_128 = cellUnderTest_io_out_ready & cellUnderTest_io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_129 = _T_127 & _T_128; // @[CFARCoreWithASR.scala 170:40]
  assign maybeFullLead_0 = _T_108; // @[CFARCoreWithASR.scala 132:32]
  assign _T_130 = leadWindow_io_regFull | maybeFullLead_0; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_739 = {{4{leadWindow_io_in_bits[15]}},leadWindow_io_in_bits}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_133 = $signed(sumSubLeads_0) + $signed(_GEN_739); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_740 = {{4{minusOperandLead[15]}},minusOperandLead}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_136 = $signed(_T_133) - $signed(_GEN_740); // @[FixedPointTypeClass.scala 30:68]
  assign _T_141 = 7'h3 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex = _T_141 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_145 = endIndex <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_146 = _T_86 & _T_145; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_1 = _T_86 ? $signed(laggWindow_io_parallelOut_7) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_1 = _T_86 ? $signed(leadWindow_io_parallelOut_7) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_148 = endIndex - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_149 = leadWindow_io_cnt > _T_148; // @[CFARCoreWithASR.scala 132:57]
  assign _T_152 = laggWindow_io_cnt > _T_148; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_1 = _T_152; // @[CFARCoreWithASR.scala 133:32]
  assign _T_156 = laggWindow_io_regFull | maybeFullLagg_1; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_742 = {{4{laggWindow_io_parallelOut_3[15]}},laggWindow_io_parallelOut_3}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_159 = $signed(sumSubLaggs_1) + $signed(_GEN_742); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_743 = {{4{minusOperandLagg_1[15]}},minusOperandLagg_1}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_162 = $signed(_T_159) - $signed(_GEN_743); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_1 = _T_149; // @[CFARCoreWithASR.scala 132:32]
  assign _T_171 = leadWindow_io_regFull | maybeFullLead_1; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_745 = {{4{leadWindow_io_parallelOut_3[15]}},leadWindow_io_parallelOut_3}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_174 = $signed(sumSubLeads_1) + $signed(_GEN_745); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_746 = {{4{minusOperandLead_1[15]}},minusOperandLead_1}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_177 = $signed(_T_174) - $signed(_GEN_746); // @[FixedPointTypeClass.scala 30:68]
  assign _T_182 = 7'h7 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_1 = _T_182 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_188 = endIndex_1 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_189 = _T_92 & _T_188; // @[CFARCoreWithASR.scala 110:64]
  assign _T_190 = _T_87 ? $signed(laggWindow_io_parallelOut_15) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLagg_2 = _T_86 ? $signed(laggWindow_io_parallelOut_11) : $signed(_T_190); // @[Mux.scala 87:16]
  assign _T_191 = _T_87 ? $signed(leadWindow_io_parallelOut_15) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_2 = _T_86 ? $signed(leadWindow_io_parallelOut_11) : $signed(_T_191); // @[Mux.scala 87:16]
  assign _T_193 = endIndex_1 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_194 = leadWindow_io_cnt > _T_193; // @[CFARCoreWithASR.scala 132:57]
  assign _T_197 = laggWindow_io_cnt > _T_193; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_2 = _T_197; // @[CFARCoreWithASR.scala 133:32]
  assign _T_201 = laggWindow_io_regFull | maybeFullLagg_2; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_748 = {{4{laggWindow_io_parallelOut_7[15]}},laggWindow_io_parallelOut_7}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_204 = $signed(sumSubLaggs_2) + $signed(_GEN_748); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_749 = {{4{minusOperandLagg_2[15]}},minusOperandLagg_2}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_207 = $signed(_T_204) - $signed(_GEN_749); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_2 = _T_194; // @[CFARCoreWithASR.scala 132:32]
  assign _T_216 = leadWindow_io_regFull | maybeFullLead_2; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_751 = {{4{leadWindow_io_parallelOut_7[15]}},leadWindow_io_parallelOut_7}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_219 = $signed(sumSubLeads_2) + $signed(_GEN_751); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_752 = {{4{minusOperandLead_2[15]}},minusOperandLead_2}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_222 = $signed(_T_219) - $signed(_GEN_752); // @[FixedPointTypeClass.scala 30:68]
  assign _T_227 = 7'hb + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_2 = _T_227 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_231 = endIndex_2 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_232 = _T_86 & _T_231; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_3 = _T_86 ? $signed(laggWindow_io_parallelOut_15) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_3 = _T_86 ? $signed(leadWindow_io_parallelOut_15) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_234 = endIndex_2 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_235 = leadWindow_io_cnt > _T_234; // @[CFARCoreWithASR.scala 132:57]
  assign _T_238 = laggWindow_io_cnt > _T_234; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_3 = _T_238; // @[CFARCoreWithASR.scala 133:32]
  assign _T_242 = laggWindow_io_regFull | maybeFullLagg_3; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_754 = {{4{laggWindow_io_parallelOut_11[15]}},laggWindow_io_parallelOut_11}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_245 = $signed(sumSubLaggs_3) + $signed(_GEN_754); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_755 = {{4{minusOperandLagg_3[15]}},minusOperandLagg_3}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_248 = $signed(_T_245) - $signed(_GEN_755); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_3 = _T_235; // @[CFARCoreWithASR.scala 132:32]
  assign _T_257 = leadWindow_io_regFull | maybeFullLead_3; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_757 = {{4{leadWindow_io_parallelOut_11[15]}},leadWindow_io_parallelOut_11}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_260 = $signed(sumSubLeads_3) + $signed(_GEN_757); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_758 = {{4{minusOperandLead_3[15]}},minusOperandLead_3}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_263 = $signed(_T_260) - $signed(_GEN_758); // @[FixedPointTypeClass.scala 30:68]
  assign _T_268 = 7'hf + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_3 = _T_268 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_276 = endIndex_3 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_277 = _T_93 & _T_276; // @[CFARCoreWithASR.scala 110:64]
  assign _T_278 = _T_88 ? $signed(laggWindow_io_parallelOut_31) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_279 = _T_87 ? $signed(laggWindow_io_parallelOut_23) : $signed(_T_278); // @[Mux.scala 87:16]
  assign minusOperandLagg_4 = _T_86 ? $signed(laggWindow_io_parallelOut_19) : $signed(_T_279); // @[Mux.scala 87:16]
  assign _T_280 = _T_88 ? $signed(leadWindow_io_parallelOut_31) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_281 = _T_87 ? $signed(leadWindow_io_parallelOut_23) : $signed(_T_280); // @[Mux.scala 87:16]
  assign minusOperandLead_4 = _T_86 ? $signed(leadWindow_io_parallelOut_19) : $signed(_T_281); // @[Mux.scala 87:16]
  assign _T_283 = endIndex_3 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_284 = leadWindow_io_cnt > _T_283; // @[CFARCoreWithASR.scala 132:57]
  assign _T_287 = laggWindow_io_cnt > _T_283; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_4 = _T_287; // @[CFARCoreWithASR.scala 133:32]
  assign _T_291 = laggWindow_io_regFull | maybeFullLagg_4; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_760 = {{4{laggWindow_io_parallelOut_15[15]}},laggWindow_io_parallelOut_15}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_294 = $signed(sumSubLaggs_4) + $signed(_GEN_760); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_761 = {{4{minusOperandLagg_4[15]}},minusOperandLagg_4}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_297 = $signed(_T_294) - $signed(_GEN_761); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_4 = _T_284; // @[CFARCoreWithASR.scala 132:32]
  assign _T_306 = leadWindow_io_regFull | maybeFullLead_4; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_763 = {{4{leadWindow_io_parallelOut_15[15]}},leadWindow_io_parallelOut_15}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_309 = $signed(sumSubLeads_4) + $signed(_GEN_763); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_764 = {{4{minusOperandLead_4[15]}},minusOperandLead_4}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_312 = $signed(_T_309) - $signed(_GEN_764); // @[FixedPointTypeClass.scala 30:68]
  assign _T_317 = 7'h13 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_4 = _T_317 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_321 = endIndex_4 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_322 = _T_86 & _T_321; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_5 = _T_86 ? $signed(laggWindow_io_parallelOut_23) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_5 = _T_86 ? $signed(leadWindow_io_parallelOut_23) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_324 = endIndex_4 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_325 = leadWindow_io_cnt > _T_324; // @[CFARCoreWithASR.scala 132:57]
  assign _T_328 = laggWindow_io_cnt > _T_324; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_5 = _T_328; // @[CFARCoreWithASR.scala 133:32]
  assign _T_332 = laggWindow_io_regFull | maybeFullLagg_5; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_766 = {{4{laggWindow_io_parallelOut_19[15]}},laggWindow_io_parallelOut_19}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_335 = $signed(sumSubLaggs_5) + $signed(_GEN_766); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_767 = {{4{minusOperandLagg_5[15]}},minusOperandLagg_5}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_338 = $signed(_T_335) - $signed(_GEN_767); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_5 = _T_325; // @[CFARCoreWithASR.scala 132:32]
  assign _T_347 = leadWindow_io_regFull | maybeFullLead_5; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_769 = {{4{leadWindow_io_parallelOut_19[15]}},leadWindow_io_parallelOut_19}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_350 = $signed(sumSubLeads_5) + $signed(_GEN_769); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_770 = {{4{minusOperandLead_5[15]}},minusOperandLead_5}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_353 = $signed(_T_350) - $signed(_GEN_770); // @[FixedPointTypeClass.scala 30:68]
  assign _T_358 = 7'h17 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_5 = _T_358 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_364 = endIndex_5 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_365 = _T_92 & _T_364; // @[CFARCoreWithASR.scala 110:64]
  assign _T_366 = _T_87 ? $signed(laggWindow_io_parallelOut_31) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLagg_6 = _T_86 ? $signed(laggWindow_io_parallelOut_27) : $signed(_T_366); // @[Mux.scala 87:16]
  assign _T_367 = _T_87 ? $signed(leadWindow_io_parallelOut_31) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_6 = _T_86 ? $signed(leadWindow_io_parallelOut_27) : $signed(_T_367); // @[Mux.scala 87:16]
  assign _T_369 = endIndex_5 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_370 = leadWindow_io_cnt > _T_369; // @[CFARCoreWithASR.scala 132:57]
  assign _T_373 = laggWindow_io_cnt > _T_369; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_6 = _T_373; // @[CFARCoreWithASR.scala 133:32]
  assign _T_377 = laggWindow_io_regFull | maybeFullLagg_6; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_772 = {{4{laggWindow_io_parallelOut_23[15]}},laggWindow_io_parallelOut_23}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_380 = $signed(sumSubLaggs_6) + $signed(_GEN_772); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_773 = {{4{minusOperandLagg_6[15]}},minusOperandLagg_6}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_383 = $signed(_T_380) - $signed(_GEN_773); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_6 = _T_370; // @[CFARCoreWithASR.scala 132:32]
  assign _T_392 = leadWindow_io_regFull | maybeFullLead_6; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_775 = {{4{leadWindow_io_parallelOut_23[15]}},leadWindow_io_parallelOut_23}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_395 = $signed(sumSubLeads_6) + $signed(_GEN_775); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_776 = {{4{minusOperandLead_6[15]}},minusOperandLead_6}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_398 = $signed(_T_395) - $signed(_GEN_776); // @[FixedPointTypeClass.scala 30:68]
  assign _T_403 = 7'h1b + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_6 = _T_403 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_407 = endIndex_6 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_408 = _T_86 & _T_407; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_7 = _T_86 ? $signed(laggWindow_io_parallelOut_31) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_7 = _T_86 ? $signed(leadWindow_io_parallelOut_31) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_410 = endIndex_6 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_411 = leadWindow_io_cnt > _T_410; // @[CFARCoreWithASR.scala 132:57]
  assign _T_414 = laggWindow_io_cnt > _T_410; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_7 = _T_414; // @[CFARCoreWithASR.scala 133:32]
  assign _T_418 = laggWindow_io_regFull | maybeFullLagg_7; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_778 = {{4{laggWindow_io_parallelOut_27[15]}},laggWindow_io_parallelOut_27}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_421 = $signed(sumSubLaggs_7) + $signed(_GEN_778); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_779 = {{4{minusOperandLagg_7[15]}},minusOperandLagg_7}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_424 = $signed(_T_421) - $signed(_GEN_779); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_7 = _T_411; // @[CFARCoreWithASR.scala 132:32]
  assign _T_433 = leadWindow_io_regFull | maybeFullLead_7; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_781 = {{4{leadWindow_io_parallelOut_27[15]}},leadWindow_io_parallelOut_27}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_436 = $signed(sumSubLeads_7) + $signed(_GEN_781); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_782 = {{4{minusOperandLead_7[15]}},minusOperandLead_7}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_439 = $signed(_T_436) - $signed(_GEN_782); // @[FixedPointTypeClass.scala 30:68]
  assign _T_444 = 7'h1f + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_7 = _T_444 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_454 = endIndex_7 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_455 = _T_94 & _T_454; // @[CFARCoreWithASR.scala 110:64]
  assign _T_456 = _T_89 ? $signed(laggWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_457 = _T_88 ? $signed(laggWindow_io_parallelOut_47) : $signed(_T_456); // @[Mux.scala 87:16]
  assign _T_458 = _T_87 ? $signed(laggWindow_io_parallelOut_39) : $signed(_T_457); // @[Mux.scala 87:16]
  assign minusOperandLagg_8 = _T_86 ? $signed(laggWindow_io_parallelOut_35) : $signed(_T_458); // @[Mux.scala 87:16]
  assign _T_459 = _T_89 ? $signed(leadWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_460 = _T_88 ? $signed(leadWindow_io_parallelOut_47) : $signed(_T_459); // @[Mux.scala 87:16]
  assign _T_461 = _T_87 ? $signed(leadWindow_io_parallelOut_39) : $signed(_T_460); // @[Mux.scala 87:16]
  assign minusOperandLead_8 = _T_86 ? $signed(leadWindow_io_parallelOut_35) : $signed(_T_461); // @[Mux.scala 87:16]
  assign _T_463 = endIndex_7 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_464 = leadWindow_io_cnt > _T_463; // @[CFARCoreWithASR.scala 132:57]
  assign _T_467 = laggWindow_io_cnt > _T_463; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_8 = _T_467; // @[CFARCoreWithASR.scala 133:32]
  assign _T_471 = laggWindow_io_regFull | maybeFullLagg_8; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_784 = {{4{laggWindow_io_parallelOut_31[15]}},laggWindow_io_parallelOut_31}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_474 = $signed(sumSubLaggs_8) + $signed(_GEN_784); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_785 = {{4{minusOperandLagg_8[15]}},minusOperandLagg_8}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_477 = $signed(_T_474) - $signed(_GEN_785); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_8 = _T_464; // @[CFARCoreWithASR.scala 132:32]
  assign _T_486 = leadWindow_io_regFull | maybeFullLead_8; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_787 = {{4{leadWindow_io_parallelOut_31[15]}},leadWindow_io_parallelOut_31}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_489 = $signed(sumSubLeads_8) + $signed(_GEN_787); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_788 = {{4{minusOperandLead_8[15]}},minusOperandLead_8}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_492 = $signed(_T_489) - $signed(_GEN_788); // @[FixedPointTypeClass.scala 30:68]
  assign _T_497 = 7'h23 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_8 = _T_497 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_501 = endIndex_8 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_502 = _T_86 & _T_501; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_9 = _T_86 ? $signed(laggWindow_io_parallelOut_39) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_9 = _T_86 ? $signed(leadWindow_io_parallelOut_39) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_504 = endIndex_8 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_505 = leadWindow_io_cnt > _T_504; // @[CFARCoreWithASR.scala 132:57]
  assign _T_508 = laggWindow_io_cnt > _T_504; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_9 = _T_508; // @[CFARCoreWithASR.scala 133:32]
  assign _T_512 = laggWindow_io_regFull | maybeFullLagg_9; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_790 = {{4{laggWindow_io_parallelOut_35[15]}},laggWindow_io_parallelOut_35}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_515 = $signed(sumSubLaggs_9) + $signed(_GEN_790); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_791 = {{4{minusOperandLagg_9[15]}},minusOperandLagg_9}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_518 = $signed(_T_515) - $signed(_GEN_791); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_9 = _T_505; // @[CFARCoreWithASR.scala 132:32]
  assign _T_527 = leadWindow_io_regFull | maybeFullLead_9; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_793 = {{4{leadWindow_io_parallelOut_35[15]}},leadWindow_io_parallelOut_35}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_530 = $signed(sumSubLeads_9) + $signed(_GEN_793); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_794 = {{4{minusOperandLead_9[15]}},minusOperandLead_9}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_533 = $signed(_T_530) - $signed(_GEN_794); // @[FixedPointTypeClass.scala 30:68]
  assign _T_538 = 7'h27 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_9 = _T_538 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_544 = endIndex_9 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_545 = _T_92 & _T_544; // @[CFARCoreWithASR.scala 110:64]
  assign _T_546 = _T_87 ? $signed(laggWindow_io_parallelOut_47) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLagg_10 = _T_86 ? $signed(laggWindow_io_parallelOut_43) : $signed(_T_546); // @[Mux.scala 87:16]
  assign _T_547 = _T_87 ? $signed(leadWindow_io_parallelOut_47) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_10 = _T_86 ? $signed(leadWindow_io_parallelOut_43) : $signed(_T_547); // @[Mux.scala 87:16]
  assign _T_549 = endIndex_9 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_550 = leadWindow_io_cnt > _T_549; // @[CFARCoreWithASR.scala 132:57]
  assign _T_553 = laggWindow_io_cnt > _T_549; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_10 = _T_553; // @[CFARCoreWithASR.scala 133:32]
  assign _T_557 = laggWindow_io_regFull | maybeFullLagg_10; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_796 = {{4{laggWindow_io_parallelOut_39[15]}},laggWindow_io_parallelOut_39}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_560 = $signed(sumSubLaggs_10) + $signed(_GEN_796); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_797 = {{4{minusOperandLagg_10[15]}},minusOperandLagg_10}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_563 = $signed(_T_560) - $signed(_GEN_797); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_10 = _T_550; // @[CFARCoreWithASR.scala 132:32]
  assign _T_572 = leadWindow_io_regFull | maybeFullLead_10; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_799 = {{4{leadWindow_io_parallelOut_39[15]}},leadWindow_io_parallelOut_39}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_575 = $signed(sumSubLeads_10) + $signed(_GEN_799); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_800 = {{4{minusOperandLead_10[15]}},minusOperandLead_10}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_578 = $signed(_T_575) - $signed(_GEN_800); // @[FixedPointTypeClass.scala 30:68]
  assign _T_583 = 7'h2b + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_10 = _T_583 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_587 = endIndex_10 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_588 = _T_86 & _T_587; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_11 = _T_86 ? $signed(laggWindow_io_parallelOut_47) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_11 = _T_86 ? $signed(leadWindow_io_parallelOut_47) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_590 = endIndex_10 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_591 = leadWindow_io_cnt > _T_590; // @[CFARCoreWithASR.scala 132:57]
  assign _T_594 = laggWindow_io_cnt > _T_590; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_11 = _T_594; // @[CFARCoreWithASR.scala 133:32]
  assign _T_598 = laggWindow_io_regFull | maybeFullLagg_11; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_802 = {{4{laggWindow_io_parallelOut_43[15]}},laggWindow_io_parallelOut_43}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_601 = $signed(sumSubLaggs_11) + $signed(_GEN_802); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_803 = {{4{minusOperandLagg_11[15]}},minusOperandLagg_11}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_604 = $signed(_T_601) - $signed(_GEN_803); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_11 = _T_591; // @[CFARCoreWithASR.scala 132:32]
  assign _T_613 = leadWindow_io_regFull | maybeFullLead_11; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_805 = {{4{leadWindow_io_parallelOut_43[15]}},leadWindow_io_parallelOut_43}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_616 = $signed(sumSubLeads_11) + $signed(_GEN_805); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_806 = {{4{minusOperandLead_11[15]}},minusOperandLead_11}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_619 = $signed(_T_616) - $signed(_GEN_806); // @[FixedPointTypeClass.scala 30:68]
  assign _T_624 = 7'h2f + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_11 = _T_624 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_632 = endIndex_11 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_633 = _T_93 & _T_632; // @[CFARCoreWithASR.scala 110:64]
  assign _T_634 = _T_88 ? $signed(laggWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_635 = _T_87 ? $signed(laggWindow_io_parallelOut_55) : $signed(_T_634); // @[Mux.scala 87:16]
  assign minusOperandLagg_12 = _T_86 ? $signed(laggWindow_io_parallelOut_51) : $signed(_T_635); // @[Mux.scala 87:16]
  assign _T_636 = _T_88 ? $signed(leadWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_637 = _T_87 ? $signed(leadWindow_io_parallelOut_55) : $signed(_T_636); // @[Mux.scala 87:16]
  assign minusOperandLead_12 = _T_86 ? $signed(leadWindow_io_parallelOut_51) : $signed(_T_637); // @[Mux.scala 87:16]
  assign _T_639 = endIndex_11 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_640 = leadWindow_io_cnt > _T_639; // @[CFARCoreWithASR.scala 132:57]
  assign _T_643 = laggWindow_io_cnt > _T_639; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_12 = _T_643; // @[CFARCoreWithASR.scala 133:32]
  assign _T_647 = laggWindow_io_regFull | maybeFullLagg_12; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_808 = {{4{laggWindow_io_parallelOut_47[15]}},laggWindow_io_parallelOut_47}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_650 = $signed(sumSubLaggs_12) + $signed(_GEN_808); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_809 = {{4{minusOperandLagg_12[15]}},minusOperandLagg_12}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_653 = $signed(_T_650) - $signed(_GEN_809); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_12 = _T_640; // @[CFARCoreWithASR.scala 132:32]
  assign _T_662 = leadWindow_io_regFull | maybeFullLead_12; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_811 = {{4{leadWindow_io_parallelOut_47[15]}},leadWindow_io_parallelOut_47}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_665 = $signed(sumSubLeads_12) + $signed(_GEN_811); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_812 = {{4{minusOperandLead_12[15]}},minusOperandLead_12}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_668 = $signed(_T_665) - $signed(_GEN_812); // @[FixedPointTypeClass.scala 30:68]
  assign _T_673 = 7'h33 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_12 = _T_673 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_677 = endIndex_12 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_678 = _T_86 & _T_677; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_13 = _T_86 ? $signed(laggWindow_io_parallelOut_55) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_13 = _T_86 ? $signed(leadWindow_io_parallelOut_55) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_680 = endIndex_12 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_681 = leadWindow_io_cnt > _T_680; // @[CFARCoreWithASR.scala 132:57]
  assign _T_684 = laggWindow_io_cnt > _T_680; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_13 = _T_684; // @[CFARCoreWithASR.scala 133:32]
  assign _T_688 = laggWindow_io_regFull | maybeFullLagg_13; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_814 = {{4{laggWindow_io_parallelOut_51[15]}},laggWindow_io_parallelOut_51}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_691 = $signed(sumSubLaggs_13) + $signed(_GEN_814); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_815 = {{4{minusOperandLagg_13[15]}},minusOperandLagg_13}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_694 = $signed(_T_691) - $signed(_GEN_815); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_13 = _T_681; // @[CFARCoreWithASR.scala 132:32]
  assign _T_703 = leadWindow_io_regFull | maybeFullLead_13; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_817 = {{4{leadWindow_io_parallelOut_51[15]}},leadWindow_io_parallelOut_51}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_706 = $signed(sumSubLeads_13) + $signed(_GEN_817); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_818 = {{4{minusOperandLead_13[15]}},minusOperandLead_13}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_709 = $signed(_T_706) - $signed(_GEN_818); // @[FixedPointTypeClass.scala 30:68]
  assign _T_714 = 7'h37 + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_13 = _T_714 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_720 = endIndex_13 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_721 = _T_92 & _T_720; // @[CFARCoreWithASR.scala 110:64]
  assign _T_722 = _T_87 ? $signed(laggWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLagg_14 = _T_86 ? $signed(laggWindow_io_parallelOut_59) : $signed(_T_722); // @[Mux.scala 87:16]
  assign _T_723 = _T_87 ? $signed(leadWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_14 = _T_86 ? $signed(leadWindow_io_parallelOut_59) : $signed(_T_723); // @[Mux.scala 87:16]
  assign _T_725 = endIndex_13 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_726 = leadWindow_io_cnt > _T_725; // @[CFARCoreWithASR.scala 132:57]
  assign _T_729 = laggWindow_io_cnt > _T_725; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_14 = _T_729; // @[CFARCoreWithASR.scala 133:32]
  assign _T_733 = laggWindow_io_regFull | maybeFullLagg_14; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_820 = {{4{laggWindow_io_parallelOut_55[15]}},laggWindow_io_parallelOut_55}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_736 = $signed(sumSubLaggs_14) + $signed(_GEN_820); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_821 = {{4{minusOperandLagg_14[15]}},minusOperandLagg_14}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_739 = $signed(_T_736) - $signed(_GEN_821); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_14 = _T_726; // @[CFARCoreWithASR.scala 132:32]
  assign _T_748 = leadWindow_io_regFull | maybeFullLead_14; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_823 = {{4{leadWindow_io_parallelOut_55[15]}},leadWindow_io_parallelOut_55}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_751 = $signed(sumSubLeads_14) + $signed(_GEN_823); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_824 = {{4{minusOperandLead_14[15]}},minusOperandLead_14}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_754 = $signed(_T_751) - $signed(_GEN_824); // @[FixedPointTypeClass.scala 30:68]
  assign _T_759 = 7'h3b + io_subCells; // @[CFARCoreWithASR.scala 103:76]
  assign endIndex_14 = _T_759 + 7'h1; // @[CFARCoreWithASR.scala 103:94]
  assign _T_763 = endIndex_14 <= io_windowCells; // @[CFARCoreWithASR.scala 110:76]
  assign _T_764 = _T_86 & _T_763; // @[CFARCoreWithASR.scala 110:64]
  assign minusOperandLagg_15 = _T_86 ? $signed(laggWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign minusOperandLead_15 = _T_86 ? $signed(leadWindow_io_parallelOut_63) : $signed(16'sh0); // @[Mux.scala 87:16]
  assign _T_766 = endIndex_14 - 7'h1; // @[CFARCoreWithASR.scala 132:69]
  assign _T_767 = leadWindow_io_cnt > _T_766; // @[CFARCoreWithASR.scala 132:57]
  assign _T_770 = laggWindow_io_cnt > _T_766; // @[CFARCoreWithASR.scala 133:57]
  assign maybeFullLagg_15 = _T_770; // @[CFARCoreWithASR.scala 133:32]
  assign _T_774 = laggWindow_io_regFull | maybeFullLagg_15; // @[CFARCoreWithASR.scala 147:35]
  assign _GEN_826 = {{4{laggWindow_io_parallelOut_59[15]}},laggWindow_io_parallelOut_59}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_777 = $signed(sumSubLaggs_15) + $signed(_GEN_826); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_827 = {{4{minusOperandLagg_15[15]}},minusOperandLagg_15}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_780 = $signed(_T_777) - $signed(_GEN_827); // @[FixedPointTypeClass.scala 30:68]
  assign maybeFullLead_15 = _T_767; // @[CFARCoreWithASR.scala 132:32]
  assign _T_789 = leadWindow_io_regFull | maybeFullLead_15; // @[CFARCoreWithASR.scala 172:35]
  assign _GEN_829 = {{4{leadWindow_io_parallelOut_59[15]}},leadWindow_io_parallelOut_59}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_792 = $signed(sumSubLeads_15) + $signed(_GEN_829); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_830 = {{4{minusOperandLead_15[15]}},minusOperandLead_15}; // @[FixedPointTypeClass.scala 30:68]
  assign _T_795 = $signed(_T_792) - $signed(_GEN_830); // @[FixedPointTypeClass.scala 30:68]
  assign _T_801 = io_subCells[6:4] != 3'h0; // @[CircuitMath.scala 37:22]
  assign _T_804 = io_subCells[6] ? 2'h2 : {{1'd0}, io_subCells[5]}; // @[CircuitMath.scala 32:10]
  assign _T_808 = io_subCells[2] ? 2'h2 : {{1'd0}, io_subCells[1]}; // @[CircuitMath.scala 32:10]
  assign _T_809 = io_subCells[3] ? 2'h3 : _T_808; // @[CircuitMath.scala 32:10]
  assign _T_810 = _T_801 ? _T_804 : _T_809; // @[CircuitMath.scala 38:21]
  assign _T_811 = {_T_801,_T_810}; // @[Cat.scala 29:58]
  assign diffInSubSize = _T_811 - 3'h2; // @[CFARCoreWithASR.scala 193:45]
  assign _T_814 = $signed(sumSubLaggs_0) > $signed(sumSubLeads_0); // @[FixedPointTypeClass.scala 55:59]
  assign max_0 = _T_814 ? $signed(sumSubLaggs_0) : $signed(sumSubLeads_0); // @[Order.scala 56:31]
  assign _T_815 = $signed(sumSubLaggs_1) > $signed(sumSubLeads_1); // @[FixedPointTypeClass.scala 55:59]
  assign max_1 = _T_815 ? $signed(sumSubLaggs_1) : $signed(sumSubLeads_1); // @[Order.scala 56:31]
  assign _T_816 = $signed(sumSubLaggs_2) > $signed(sumSubLeads_2); // @[FixedPointTypeClass.scala 55:59]
  assign max_2 = _T_816 ? $signed(sumSubLaggs_2) : $signed(sumSubLeads_2); // @[Order.scala 56:31]
  assign _T_817 = $signed(sumSubLaggs_3) > $signed(sumSubLeads_3); // @[FixedPointTypeClass.scala 55:59]
  assign max_3 = _T_817 ? $signed(sumSubLaggs_3) : $signed(sumSubLeads_3); // @[Order.scala 56:31]
  assign _T_818 = $signed(sumSubLaggs_4) > $signed(sumSubLeads_4); // @[FixedPointTypeClass.scala 55:59]
  assign max_4 = _T_818 ? $signed(sumSubLaggs_4) : $signed(sumSubLeads_4); // @[Order.scala 56:31]
  assign _T_819 = $signed(sumSubLaggs_5) > $signed(sumSubLeads_5); // @[FixedPointTypeClass.scala 55:59]
  assign max_5 = _T_819 ? $signed(sumSubLaggs_5) : $signed(sumSubLeads_5); // @[Order.scala 56:31]
  assign _T_820 = $signed(sumSubLaggs_6) > $signed(sumSubLeads_6); // @[FixedPointTypeClass.scala 55:59]
  assign max_6 = _T_820 ? $signed(sumSubLaggs_6) : $signed(sumSubLeads_6); // @[Order.scala 56:31]
  assign _T_821 = $signed(sumSubLaggs_7) > $signed(sumSubLeads_7); // @[FixedPointTypeClass.scala 55:59]
  assign max_7 = _T_821 ? $signed(sumSubLaggs_7) : $signed(sumSubLeads_7); // @[Order.scala 56:31]
  assign _T_822 = $signed(sumSubLaggs_8) > $signed(sumSubLeads_8); // @[FixedPointTypeClass.scala 55:59]
  assign max_8 = _T_822 ? $signed(sumSubLaggs_8) : $signed(sumSubLeads_8); // @[Order.scala 56:31]
  assign _T_823 = $signed(sumSubLaggs_9) > $signed(sumSubLeads_9); // @[FixedPointTypeClass.scala 55:59]
  assign max_9 = _T_823 ? $signed(sumSubLaggs_9) : $signed(sumSubLeads_9); // @[Order.scala 56:31]
  assign _T_824 = $signed(sumSubLaggs_10) > $signed(sumSubLeads_10); // @[FixedPointTypeClass.scala 55:59]
  assign max_10 = _T_824 ? $signed(sumSubLaggs_10) : $signed(sumSubLeads_10); // @[Order.scala 56:31]
  assign _T_825 = $signed(sumSubLaggs_11) > $signed(sumSubLeads_11); // @[FixedPointTypeClass.scala 55:59]
  assign max_11 = _T_825 ? $signed(sumSubLaggs_11) : $signed(sumSubLeads_11); // @[Order.scala 56:31]
  assign _T_826 = $signed(sumSubLaggs_12) > $signed(sumSubLeads_12); // @[FixedPointTypeClass.scala 55:59]
  assign max_12 = _T_826 ? $signed(sumSubLaggs_12) : $signed(sumSubLeads_12); // @[Order.scala 56:31]
  assign _T_827 = $signed(sumSubLaggs_13) > $signed(sumSubLeads_13); // @[FixedPointTypeClass.scala 55:59]
  assign max_13 = _T_827 ? $signed(sumSubLaggs_13) : $signed(sumSubLeads_13); // @[Order.scala 56:31]
  assign _T_828 = $signed(sumSubLaggs_14) > $signed(sumSubLeads_14); // @[FixedPointTypeClass.scala 55:59]
  assign max_14 = _T_828 ? $signed(sumSubLaggs_14) : $signed(sumSubLeads_14); // @[Order.scala 56:31]
  assign _T_829 = $signed(sumSubLaggs_15) > $signed(sumSubLeads_15); // @[FixedPointTypeClass.scala 55:59]
  assign max_15 = _T_829 ? $signed(sumSubLaggs_15) : $signed(sumSubLeads_15); // @[Order.scala 56:31]
  assign activeSums_0 = _T_97; // @[CFARCoreWithASR.scala 110:29]
  assign _T_864 = 1'h0 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_127 = ~_T_864 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_128 = _T_864 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_832 = {{1'd0}, _T_864}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_129 = 2'h2 == _GEN_832 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_130 = 2'h3 == _GEN_832 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_834 = {{2'd0}, _T_864}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_131 = 3'h4 == _GEN_834 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_132 = 3'h5 == _GEN_834 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_133 = 3'h6 == _GEN_834 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_134 = 3'h7 == _GEN_834 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_838 = {{3'd0}, _T_864}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_135 = 4'h8 == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_136 = 4'h9 == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_137 = 4'ha == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_138 = 4'hb == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_139 = 4'hc == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_140 = 4'hd == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_141 = 4'he == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_142 = 4'hf == _GEN_838 ? $signed(max_0) : $signed(20'sh0); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_143 = activeSums_0 ? $signed(_GEN_127) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_144 = activeSums_0 ? $signed(_GEN_128) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_145 = activeSums_0 ? $signed(_GEN_129) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_146 = activeSums_0 ? $signed(_GEN_130) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_147 = activeSums_0 ? $signed(_GEN_131) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_148 = activeSums_0 ? $signed(_GEN_132) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_149 = activeSums_0 ? $signed(_GEN_133) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_150 = activeSums_0 ? $signed(_GEN_134) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_151 = activeSums_0 ? $signed(_GEN_135) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_152 = activeSums_0 ? $signed(_GEN_136) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_153 = activeSums_0 ? $signed(_GEN_137) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_154 = activeSums_0 ? $signed(_GEN_138) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_155 = activeSums_0 ? $signed(_GEN_139) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_156 = activeSums_0 ? $signed(_GEN_140) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_157 = activeSums_0 ? $signed(_GEN_141) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_158 = activeSums_0 ? $signed(_GEN_142) : $signed(20'sh0); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_1 = _T_146; // @[CFARCoreWithASR.scala 110:29]
  assign _T_866 = 1'h1 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_159 = ~_T_866 ? $signed(max_1) : $signed(_GEN_143); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_160 = _T_866 ? $signed(max_1) : $signed(_GEN_144); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_846 = {{1'd0}, _T_866}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_161 = 2'h2 == _GEN_846 ? $signed(max_1) : $signed(_GEN_145); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_162 = 2'h3 == _GEN_846 ? $signed(max_1) : $signed(_GEN_146); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_848 = {{2'd0}, _T_866}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_163 = 3'h4 == _GEN_848 ? $signed(max_1) : $signed(_GEN_147); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_164 = 3'h5 == _GEN_848 ? $signed(max_1) : $signed(_GEN_148); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_165 = 3'h6 == _GEN_848 ? $signed(max_1) : $signed(_GEN_149); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_166 = 3'h7 == _GEN_848 ? $signed(max_1) : $signed(_GEN_150); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_852 = {{3'd0}, _T_866}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_167 = 4'h8 == _GEN_852 ? $signed(max_1) : $signed(_GEN_151); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_168 = 4'h9 == _GEN_852 ? $signed(max_1) : $signed(_GEN_152); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_169 = 4'ha == _GEN_852 ? $signed(max_1) : $signed(_GEN_153); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_170 = 4'hb == _GEN_852 ? $signed(max_1) : $signed(_GEN_154); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_171 = 4'hc == _GEN_852 ? $signed(max_1) : $signed(_GEN_155); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_172 = 4'hd == _GEN_852 ? $signed(max_1) : $signed(_GEN_156); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_173 = 4'he == _GEN_852 ? $signed(max_1) : $signed(_GEN_157); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_174 = 4'hf == _GEN_852 ? $signed(max_1) : $signed(_GEN_158); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_175 = activeSums_1 ? $signed(_GEN_159) : $signed(_GEN_143); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_176 = activeSums_1 ? $signed(_GEN_160) : $signed(_GEN_144); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_177 = activeSums_1 ? $signed(_GEN_161) : $signed(_GEN_145); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_178 = activeSums_1 ? $signed(_GEN_162) : $signed(_GEN_146); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_179 = activeSums_1 ? $signed(_GEN_163) : $signed(_GEN_147); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_180 = activeSums_1 ? $signed(_GEN_164) : $signed(_GEN_148); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_181 = activeSums_1 ? $signed(_GEN_165) : $signed(_GEN_149); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_182 = activeSums_1 ? $signed(_GEN_166) : $signed(_GEN_150); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_183 = activeSums_1 ? $signed(_GEN_167) : $signed(_GEN_151); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_184 = activeSums_1 ? $signed(_GEN_168) : $signed(_GEN_152); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_185 = activeSums_1 ? $signed(_GEN_169) : $signed(_GEN_153); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_186 = activeSums_1 ? $signed(_GEN_170) : $signed(_GEN_154); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_187 = activeSums_1 ? $signed(_GEN_171) : $signed(_GEN_155); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_188 = activeSums_1 ? $signed(_GEN_172) : $signed(_GEN_156); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_189 = activeSums_1 ? $signed(_GEN_173) : $signed(_GEN_157); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_190 = activeSums_1 ? $signed(_GEN_174) : $signed(_GEN_158); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_2 = _T_189; // @[CFARCoreWithASR.scala 110:29]
  assign _T_868 = 2'h2 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_191 = 2'h0 == _T_868 ? $signed(max_2) : $signed(_GEN_175); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_192 = 2'h1 == _T_868 ? $signed(max_2) : $signed(_GEN_176); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_193 = 2'h2 == _T_868 ? $signed(max_2) : $signed(_GEN_177); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_194 = 2'h3 == _T_868 ? $signed(max_2) : $signed(_GEN_178); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_860 = {{1'd0}, _T_868}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_195 = 3'h4 == _GEN_860 ? $signed(max_2) : $signed(_GEN_179); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_196 = 3'h5 == _GEN_860 ? $signed(max_2) : $signed(_GEN_180); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_197 = 3'h6 == _GEN_860 ? $signed(max_2) : $signed(_GEN_181); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_198 = 3'h7 == _GEN_860 ? $signed(max_2) : $signed(_GEN_182); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_864 = {{2'd0}, _T_868}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_199 = 4'h8 == _GEN_864 ? $signed(max_2) : $signed(_GEN_183); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_200 = 4'h9 == _GEN_864 ? $signed(max_2) : $signed(_GEN_184); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_201 = 4'ha == _GEN_864 ? $signed(max_2) : $signed(_GEN_185); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_202 = 4'hb == _GEN_864 ? $signed(max_2) : $signed(_GEN_186); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_203 = 4'hc == _GEN_864 ? $signed(max_2) : $signed(_GEN_187); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_204 = 4'hd == _GEN_864 ? $signed(max_2) : $signed(_GEN_188); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_205 = 4'he == _GEN_864 ? $signed(max_2) : $signed(_GEN_189); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_206 = 4'hf == _GEN_864 ? $signed(max_2) : $signed(_GEN_190); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_207 = activeSums_2 ? $signed(_GEN_191) : $signed(_GEN_175); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_208 = activeSums_2 ? $signed(_GEN_192) : $signed(_GEN_176); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_209 = activeSums_2 ? $signed(_GEN_193) : $signed(_GEN_177); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_210 = activeSums_2 ? $signed(_GEN_194) : $signed(_GEN_178); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_211 = activeSums_2 ? $signed(_GEN_195) : $signed(_GEN_179); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_212 = activeSums_2 ? $signed(_GEN_196) : $signed(_GEN_180); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_213 = activeSums_2 ? $signed(_GEN_197) : $signed(_GEN_181); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_214 = activeSums_2 ? $signed(_GEN_198) : $signed(_GEN_182); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_215 = activeSums_2 ? $signed(_GEN_199) : $signed(_GEN_183); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_216 = activeSums_2 ? $signed(_GEN_200) : $signed(_GEN_184); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_217 = activeSums_2 ? $signed(_GEN_201) : $signed(_GEN_185); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_218 = activeSums_2 ? $signed(_GEN_202) : $signed(_GEN_186); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_219 = activeSums_2 ? $signed(_GEN_203) : $signed(_GEN_187); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_220 = activeSums_2 ? $signed(_GEN_204) : $signed(_GEN_188); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_221 = activeSums_2 ? $signed(_GEN_205) : $signed(_GEN_189); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_222 = activeSums_2 ? $signed(_GEN_206) : $signed(_GEN_190); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_3 = _T_232; // @[CFARCoreWithASR.scala 110:29]
  assign _T_870 = 2'h3 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_223 = 2'h0 == _T_870 ? $signed(max_3) : $signed(_GEN_207); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_224 = 2'h1 == _T_870 ? $signed(max_3) : $signed(_GEN_208); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_225 = 2'h2 == _T_870 ? $signed(max_3) : $signed(_GEN_209); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_226 = 2'h3 == _T_870 ? $signed(max_3) : $signed(_GEN_210); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_872 = {{1'd0}, _T_870}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_227 = 3'h4 == _GEN_872 ? $signed(max_3) : $signed(_GEN_211); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_228 = 3'h5 == _GEN_872 ? $signed(max_3) : $signed(_GEN_212); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_229 = 3'h6 == _GEN_872 ? $signed(max_3) : $signed(_GEN_213); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_230 = 3'h7 == _GEN_872 ? $signed(max_3) : $signed(_GEN_214); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_876 = {{2'd0}, _T_870}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_231 = 4'h8 == _GEN_876 ? $signed(max_3) : $signed(_GEN_215); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_232 = 4'h9 == _GEN_876 ? $signed(max_3) : $signed(_GEN_216); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_233 = 4'ha == _GEN_876 ? $signed(max_3) : $signed(_GEN_217); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_234 = 4'hb == _GEN_876 ? $signed(max_3) : $signed(_GEN_218); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_235 = 4'hc == _GEN_876 ? $signed(max_3) : $signed(_GEN_219); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_236 = 4'hd == _GEN_876 ? $signed(max_3) : $signed(_GEN_220); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_237 = 4'he == _GEN_876 ? $signed(max_3) : $signed(_GEN_221); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_238 = 4'hf == _GEN_876 ? $signed(max_3) : $signed(_GEN_222); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_239 = activeSums_3 ? $signed(_GEN_223) : $signed(_GEN_207); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_240 = activeSums_3 ? $signed(_GEN_224) : $signed(_GEN_208); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_241 = activeSums_3 ? $signed(_GEN_225) : $signed(_GEN_209); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_242 = activeSums_3 ? $signed(_GEN_226) : $signed(_GEN_210); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_243 = activeSums_3 ? $signed(_GEN_227) : $signed(_GEN_211); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_244 = activeSums_3 ? $signed(_GEN_228) : $signed(_GEN_212); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_245 = activeSums_3 ? $signed(_GEN_229) : $signed(_GEN_213); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_246 = activeSums_3 ? $signed(_GEN_230) : $signed(_GEN_214); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_247 = activeSums_3 ? $signed(_GEN_231) : $signed(_GEN_215); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_248 = activeSums_3 ? $signed(_GEN_232) : $signed(_GEN_216); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_249 = activeSums_3 ? $signed(_GEN_233) : $signed(_GEN_217); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_250 = activeSums_3 ? $signed(_GEN_234) : $signed(_GEN_218); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_251 = activeSums_3 ? $signed(_GEN_235) : $signed(_GEN_219); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_252 = activeSums_3 ? $signed(_GEN_236) : $signed(_GEN_220); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_253 = activeSums_3 ? $signed(_GEN_237) : $signed(_GEN_221); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_254 = activeSums_3 ? $signed(_GEN_238) : $signed(_GEN_222); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_4 = _T_277; // @[CFARCoreWithASR.scala 110:29]
  assign _T_872 = 3'h4 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_255 = 3'h0 == _T_872 ? $signed(max_4) : $signed(_GEN_239); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_256 = 3'h1 == _T_872 ? $signed(max_4) : $signed(_GEN_240); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_257 = 3'h2 == _T_872 ? $signed(max_4) : $signed(_GEN_241); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_258 = 3'h3 == _T_872 ? $signed(max_4) : $signed(_GEN_242); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_259 = 3'h4 == _T_872 ? $signed(max_4) : $signed(_GEN_243); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_260 = 3'h5 == _T_872 ? $signed(max_4) : $signed(_GEN_244); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_261 = 3'h6 == _T_872 ? $signed(max_4) : $signed(_GEN_245); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_262 = 3'h7 == _T_872 ? $signed(max_4) : $signed(_GEN_246); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_884 = {{1'd0}, _T_872}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_263 = 4'h8 == _GEN_884 ? $signed(max_4) : $signed(_GEN_247); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_264 = 4'h9 == _GEN_884 ? $signed(max_4) : $signed(_GEN_248); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_265 = 4'ha == _GEN_884 ? $signed(max_4) : $signed(_GEN_249); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_266 = 4'hb == _GEN_884 ? $signed(max_4) : $signed(_GEN_250); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_267 = 4'hc == _GEN_884 ? $signed(max_4) : $signed(_GEN_251); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_268 = 4'hd == _GEN_884 ? $signed(max_4) : $signed(_GEN_252); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_269 = 4'he == _GEN_884 ? $signed(max_4) : $signed(_GEN_253); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_270 = 4'hf == _GEN_884 ? $signed(max_4) : $signed(_GEN_254); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_271 = activeSums_4 ? $signed(_GEN_255) : $signed(_GEN_239); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_272 = activeSums_4 ? $signed(_GEN_256) : $signed(_GEN_240); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_273 = activeSums_4 ? $signed(_GEN_257) : $signed(_GEN_241); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_274 = activeSums_4 ? $signed(_GEN_258) : $signed(_GEN_242); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_275 = activeSums_4 ? $signed(_GEN_259) : $signed(_GEN_243); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_276 = activeSums_4 ? $signed(_GEN_260) : $signed(_GEN_244); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_277 = activeSums_4 ? $signed(_GEN_261) : $signed(_GEN_245); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_278 = activeSums_4 ? $signed(_GEN_262) : $signed(_GEN_246); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_279 = activeSums_4 ? $signed(_GEN_263) : $signed(_GEN_247); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_280 = activeSums_4 ? $signed(_GEN_264) : $signed(_GEN_248); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_281 = activeSums_4 ? $signed(_GEN_265) : $signed(_GEN_249); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_282 = activeSums_4 ? $signed(_GEN_266) : $signed(_GEN_250); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_283 = activeSums_4 ? $signed(_GEN_267) : $signed(_GEN_251); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_284 = activeSums_4 ? $signed(_GEN_268) : $signed(_GEN_252); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_285 = activeSums_4 ? $signed(_GEN_269) : $signed(_GEN_253); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_286 = activeSums_4 ? $signed(_GEN_270) : $signed(_GEN_254); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_5 = _T_322; // @[CFARCoreWithASR.scala 110:29]
  assign _T_874 = 3'h5 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_287 = 3'h0 == _T_874 ? $signed(max_5) : $signed(_GEN_271); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_288 = 3'h1 == _T_874 ? $signed(max_5) : $signed(_GEN_272); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_289 = 3'h2 == _T_874 ? $signed(max_5) : $signed(_GEN_273); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_290 = 3'h3 == _T_874 ? $signed(max_5) : $signed(_GEN_274); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_291 = 3'h4 == _T_874 ? $signed(max_5) : $signed(_GEN_275); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_292 = 3'h5 == _T_874 ? $signed(max_5) : $signed(_GEN_276); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_293 = 3'h6 == _T_874 ? $signed(max_5) : $signed(_GEN_277); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_294 = 3'h7 == _T_874 ? $signed(max_5) : $signed(_GEN_278); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_892 = {{1'd0}, _T_874}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_295 = 4'h8 == _GEN_892 ? $signed(max_5) : $signed(_GEN_279); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_296 = 4'h9 == _GEN_892 ? $signed(max_5) : $signed(_GEN_280); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_297 = 4'ha == _GEN_892 ? $signed(max_5) : $signed(_GEN_281); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_298 = 4'hb == _GEN_892 ? $signed(max_5) : $signed(_GEN_282); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_299 = 4'hc == _GEN_892 ? $signed(max_5) : $signed(_GEN_283); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_300 = 4'hd == _GEN_892 ? $signed(max_5) : $signed(_GEN_284); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_301 = 4'he == _GEN_892 ? $signed(max_5) : $signed(_GEN_285); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_302 = 4'hf == _GEN_892 ? $signed(max_5) : $signed(_GEN_286); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_303 = activeSums_5 ? $signed(_GEN_287) : $signed(_GEN_271); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_304 = activeSums_5 ? $signed(_GEN_288) : $signed(_GEN_272); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_305 = activeSums_5 ? $signed(_GEN_289) : $signed(_GEN_273); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_306 = activeSums_5 ? $signed(_GEN_290) : $signed(_GEN_274); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_307 = activeSums_5 ? $signed(_GEN_291) : $signed(_GEN_275); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_308 = activeSums_5 ? $signed(_GEN_292) : $signed(_GEN_276); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_309 = activeSums_5 ? $signed(_GEN_293) : $signed(_GEN_277); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_310 = activeSums_5 ? $signed(_GEN_294) : $signed(_GEN_278); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_311 = activeSums_5 ? $signed(_GEN_295) : $signed(_GEN_279); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_312 = activeSums_5 ? $signed(_GEN_296) : $signed(_GEN_280); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_313 = activeSums_5 ? $signed(_GEN_297) : $signed(_GEN_281); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_314 = activeSums_5 ? $signed(_GEN_298) : $signed(_GEN_282); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_315 = activeSums_5 ? $signed(_GEN_299) : $signed(_GEN_283); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_316 = activeSums_5 ? $signed(_GEN_300) : $signed(_GEN_284); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_317 = activeSums_5 ? $signed(_GEN_301) : $signed(_GEN_285); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_318 = activeSums_5 ? $signed(_GEN_302) : $signed(_GEN_286); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_6 = _T_365; // @[CFARCoreWithASR.scala 110:29]
  assign _T_876 = 3'h6 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_319 = 3'h0 == _T_876 ? $signed(max_6) : $signed(_GEN_303); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_320 = 3'h1 == _T_876 ? $signed(max_6) : $signed(_GEN_304); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_321 = 3'h2 == _T_876 ? $signed(max_6) : $signed(_GEN_305); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_322 = 3'h3 == _T_876 ? $signed(max_6) : $signed(_GEN_306); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_323 = 3'h4 == _T_876 ? $signed(max_6) : $signed(_GEN_307); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_324 = 3'h5 == _T_876 ? $signed(max_6) : $signed(_GEN_308); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_325 = 3'h6 == _T_876 ? $signed(max_6) : $signed(_GEN_309); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_326 = 3'h7 == _T_876 ? $signed(max_6) : $signed(_GEN_310); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_900 = {{1'd0}, _T_876}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_327 = 4'h8 == _GEN_900 ? $signed(max_6) : $signed(_GEN_311); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_328 = 4'h9 == _GEN_900 ? $signed(max_6) : $signed(_GEN_312); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_329 = 4'ha == _GEN_900 ? $signed(max_6) : $signed(_GEN_313); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_330 = 4'hb == _GEN_900 ? $signed(max_6) : $signed(_GEN_314); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_331 = 4'hc == _GEN_900 ? $signed(max_6) : $signed(_GEN_315); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_332 = 4'hd == _GEN_900 ? $signed(max_6) : $signed(_GEN_316); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_333 = 4'he == _GEN_900 ? $signed(max_6) : $signed(_GEN_317); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_334 = 4'hf == _GEN_900 ? $signed(max_6) : $signed(_GEN_318); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_335 = activeSums_6 ? $signed(_GEN_319) : $signed(_GEN_303); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_336 = activeSums_6 ? $signed(_GEN_320) : $signed(_GEN_304); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_337 = activeSums_6 ? $signed(_GEN_321) : $signed(_GEN_305); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_338 = activeSums_6 ? $signed(_GEN_322) : $signed(_GEN_306); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_339 = activeSums_6 ? $signed(_GEN_323) : $signed(_GEN_307); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_340 = activeSums_6 ? $signed(_GEN_324) : $signed(_GEN_308); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_341 = activeSums_6 ? $signed(_GEN_325) : $signed(_GEN_309); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_342 = activeSums_6 ? $signed(_GEN_326) : $signed(_GEN_310); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_343 = activeSums_6 ? $signed(_GEN_327) : $signed(_GEN_311); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_344 = activeSums_6 ? $signed(_GEN_328) : $signed(_GEN_312); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_345 = activeSums_6 ? $signed(_GEN_329) : $signed(_GEN_313); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_346 = activeSums_6 ? $signed(_GEN_330) : $signed(_GEN_314); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_347 = activeSums_6 ? $signed(_GEN_331) : $signed(_GEN_315); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_348 = activeSums_6 ? $signed(_GEN_332) : $signed(_GEN_316); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_349 = activeSums_6 ? $signed(_GEN_333) : $signed(_GEN_317); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_350 = activeSums_6 ? $signed(_GEN_334) : $signed(_GEN_318); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_7 = _T_408; // @[CFARCoreWithASR.scala 110:29]
  assign _T_878 = 3'h7 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_351 = 3'h0 == _T_878 ? $signed(max_7) : $signed(_GEN_335); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_352 = 3'h1 == _T_878 ? $signed(max_7) : $signed(_GEN_336); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_353 = 3'h2 == _T_878 ? $signed(max_7) : $signed(_GEN_337); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_354 = 3'h3 == _T_878 ? $signed(max_7) : $signed(_GEN_338); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_355 = 3'h4 == _T_878 ? $signed(max_7) : $signed(_GEN_339); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_356 = 3'h5 == _T_878 ? $signed(max_7) : $signed(_GEN_340); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_357 = 3'h6 == _T_878 ? $signed(max_7) : $signed(_GEN_341); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_358 = 3'h7 == _T_878 ? $signed(max_7) : $signed(_GEN_342); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_908 = {{1'd0}, _T_878}; // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_359 = 4'h8 == _GEN_908 ? $signed(max_7) : $signed(_GEN_343); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_360 = 4'h9 == _GEN_908 ? $signed(max_7) : $signed(_GEN_344); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_361 = 4'ha == _GEN_908 ? $signed(max_7) : $signed(_GEN_345); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_362 = 4'hb == _GEN_908 ? $signed(max_7) : $signed(_GEN_346); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_363 = 4'hc == _GEN_908 ? $signed(max_7) : $signed(_GEN_347); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_364 = 4'hd == _GEN_908 ? $signed(max_7) : $signed(_GEN_348); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_365 = 4'he == _GEN_908 ? $signed(max_7) : $signed(_GEN_349); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_366 = 4'hf == _GEN_908 ? $signed(max_7) : $signed(_GEN_350); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_367 = activeSums_7 ? $signed(_GEN_351) : $signed(_GEN_335); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_368 = activeSums_7 ? $signed(_GEN_352) : $signed(_GEN_336); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_369 = activeSums_7 ? $signed(_GEN_353) : $signed(_GEN_337); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_370 = activeSums_7 ? $signed(_GEN_354) : $signed(_GEN_338); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_371 = activeSums_7 ? $signed(_GEN_355) : $signed(_GEN_339); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_372 = activeSums_7 ? $signed(_GEN_356) : $signed(_GEN_340); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_373 = activeSums_7 ? $signed(_GEN_357) : $signed(_GEN_341); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_374 = activeSums_7 ? $signed(_GEN_358) : $signed(_GEN_342); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_375 = activeSums_7 ? $signed(_GEN_359) : $signed(_GEN_343); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_376 = activeSums_7 ? $signed(_GEN_360) : $signed(_GEN_344); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_377 = activeSums_7 ? $signed(_GEN_361) : $signed(_GEN_345); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_378 = activeSums_7 ? $signed(_GEN_362) : $signed(_GEN_346); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_379 = activeSums_7 ? $signed(_GEN_363) : $signed(_GEN_347); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_380 = activeSums_7 ? $signed(_GEN_364) : $signed(_GEN_348); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_381 = activeSums_7 ? $signed(_GEN_365) : $signed(_GEN_349); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_382 = activeSums_7 ? $signed(_GEN_366) : $signed(_GEN_350); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_8 = _T_455; // @[CFARCoreWithASR.scala 110:29]
  assign _T_880 = 4'h8 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_383 = 4'h0 == _T_880 ? $signed(max_8) : $signed(_GEN_367); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_384 = 4'h1 == _T_880 ? $signed(max_8) : $signed(_GEN_368); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_385 = 4'h2 == _T_880 ? $signed(max_8) : $signed(_GEN_369); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_386 = 4'h3 == _T_880 ? $signed(max_8) : $signed(_GEN_370); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_387 = 4'h4 == _T_880 ? $signed(max_8) : $signed(_GEN_371); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_388 = 4'h5 == _T_880 ? $signed(max_8) : $signed(_GEN_372); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_389 = 4'h6 == _T_880 ? $signed(max_8) : $signed(_GEN_373); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_390 = 4'h7 == _T_880 ? $signed(max_8) : $signed(_GEN_374); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_391 = 4'h8 == _T_880 ? $signed(max_8) : $signed(_GEN_375); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_392 = 4'h9 == _T_880 ? $signed(max_8) : $signed(_GEN_376); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_393 = 4'ha == _T_880 ? $signed(max_8) : $signed(_GEN_377); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_394 = 4'hb == _T_880 ? $signed(max_8) : $signed(_GEN_378); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_395 = 4'hc == _T_880 ? $signed(max_8) : $signed(_GEN_379); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_396 = 4'hd == _T_880 ? $signed(max_8) : $signed(_GEN_380); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_397 = 4'he == _T_880 ? $signed(max_8) : $signed(_GEN_381); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_398 = 4'hf == _T_880 ? $signed(max_8) : $signed(_GEN_382); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_399 = activeSums_8 ? $signed(_GEN_383) : $signed(_GEN_367); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_400 = activeSums_8 ? $signed(_GEN_384) : $signed(_GEN_368); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_401 = activeSums_8 ? $signed(_GEN_385) : $signed(_GEN_369); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_402 = activeSums_8 ? $signed(_GEN_386) : $signed(_GEN_370); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_403 = activeSums_8 ? $signed(_GEN_387) : $signed(_GEN_371); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_404 = activeSums_8 ? $signed(_GEN_388) : $signed(_GEN_372); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_405 = activeSums_8 ? $signed(_GEN_389) : $signed(_GEN_373); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_406 = activeSums_8 ? $signed(_GEN_390) : $signed(_GEN_374); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_407 = activeSums_8 ? $signed(_GEN_391) : $signed(_GEN_375); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_408 = activeSums_8 ? $signed(_GEN_392) : $signed(_GEN_376); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_409 = activeSums_8 ? $signed(_GEN_393) : $signed(_GEN_377); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_410 = activeSums_8 ? $signed(_GEN_394) : $signed(_GEN_378); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_411 = activeSums_8 ? $signed(_GEN_395) : $signed(_GEN_379); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_412 = activeSums_8 ? $signed(_GEN_396) : $signed(_GEN_380); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_413 = activeSums_8 ? $signed(_GEN_397) : $signed(_GEN_381); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_414 = activeSums_8 ? $signed(_GEN_398) : $signed(_GEN_382); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_9 = _T_502; // @[CFARCoreWithASR.scala 110:29]
  assign _T_882 = 4'h9 >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_415 = 4'h0 == _T_882 ? $signed(max_9) : $signed(_GEN_399); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_416 = 4'h1 == _T_882 ? $signed(max_9) : $signed(_GEN_400); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_417 = 4'h2 == _T_882 ? $signed(max_9) : $signed(_GEN_401); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_418 = 4'h3 == _T_882 ? $signed(max_9) : $signed(_GEN_402); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_419 = 4'h4 == _T_882 ? $signed(max_9) : $signed(_GEN_403); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_420 = 4'h5 == _T_882 ? $signed(max_9) : $signed(_GEN_404); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_421 = 4'h6 == _T_882 ? $signed(max_9) : $signed(_GEN_405); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_422 = 4'h7 == _T_882 ? $signed(max_9) : $signed(_GEN_406); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_423 = 4'h8 == _T_882 ? $signed(max_9) : $signed(_GEN_407); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_424 = 4'h9 == _T_882 ? $signed(max_9) : $signed(_GEN_408); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_425 = 4'ha == _T_882 ? $signed(max_9) : $signed(_GEN_409); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_426 = 4'hb == _T_882 ? $signed(max_9) : $signed(_GEN_410); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_427 = 4'hc == _T_882 ? $signed(max_9) : $signed(_GEN_411); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_428 = 4'hd == _T_882 ? $signed(max_9) : $signed(_GEN_412); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_429 = 4'he == _T_882 ? $signed(max_9) : $signed(_GEN_413); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_430 = 4'hf == _T_882 ? $signed(max_9) : $signed(_GEN_414); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_431 = activeSums_9 ? $signed(_GEN_415) : $signed(_GEN_399); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_432 = activeSums_9 ? $signed(_GEN_416) : $signed(_GEN_400); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_433 = activeSums_9 ? $signed(_GEN_417) : $signed(_GEN_401); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_434 = activeSums_9 ? $signed(_GEN_418) : $signed(_GEN_402); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_435 = activeSums_9 ? $signed(_GEN_419) : $signed(_GEN_403); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_436 = activeSums_9 ? $signed(_GEN_420) : $signed(_GEN_404); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_437 = activeSums_9 ? $signed(_GEN_421) : $signed(_GEN_405); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_438 = activeSums_9 ? $signed(_GEN_422) : $signed(_GEN_406); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_439 = activeSums_9 ? $signed(_GEN_423) : $signed(_GEN_407); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_440 = activeSums_9 ? $signed(_GEN_424) : $signed(_GEN_408); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_441 = activeSums_9 ? $signed(_GEN_425) : $signed(_GEN_409); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_442 = activeSums_9 ? $signed(_GEN_426) : $signed(_GEN_410); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_443 = activeSums_9 ? $signed(_GEN_427) : $signed(_GEN_411); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_444 = activeSums_9 ? $signed(_GEN_428) : $signed(_GEN_412); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_445 = activeSums_9 ? $signed(_GEN_429) : $signed(_GEN_413); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_446 = activeSums_9 ? $signed(_GEN_430) : $signed(_GEN_414); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_10 = _T_545; // @[CFARCoreWithASR.scala 110:29]
  assign _T_884 = 4'ha >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_447 = 4'h0 == _T_884 ? $signed(max_10) : $signed(_GEN_431); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_448 = 4'h1 == _T_884 ? $signed(max_10) : $signed(_GEN_432); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_449 = 4'h2 == _T_884 ? $signed(max_10) : $signed(_GEN_433); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_450 = 4'h3 == _T_884 ? $signed(max_10) : $signed(_GEN_434); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_451 = 4'h4 == _T_884 ? $signed(max_10) : $signed(_GEN_435); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_452 = 4'h5 == _T_884 ? $signed(max_10) : $signed(_GEN_436); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_453 = 4'h6 == _T_884 ? $signed(max_10) : $signed(_GEN_437); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_454 = 4'h7 == _T_884 ? $signed(max_10) : $signed(_GEN_438); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_455 = 4'h8 == _T_884 ? $signed(max_10) : $signed(_GEN_439); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_456 = 4'h9 == _T_884 ? $signed(max_10) : $signed(_GEN_440); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_457 = 4'ha == _T_884 ? $signed(max_10) : $signed(_GEN_441); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_458 = 4'hb == _T_884 ? $signed(max_10) : $signed(_GEN_442); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_459 = 4'hc == _T_884 ? $signed(max_10) : $signed(_GEN_443); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_460 = 4'hd == _T_884 ? $signed(max_10) : $signed(_GEN_444); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_461 = 4'he == _T_884 ? $signed(max_10) : $signed(_GEN_445); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_462 = 4'hf == _T_884 ? $signed(max_10) : $signed(_GEN_446); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_463 = activeSums_10 ? $signed(_GEN_447) : $signed(_GEN_431); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_464 = activeSums_10 ? $signed(_GEN_448) : $signed(_GEN_432); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_465 = activeSums_10 ? $signed(_GEN_449) : $signed(_GEN_433); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_466 = activeSums_10 ? $signed(_GEN_450) : $signed(_GEN_434); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_467 = activeSums_10 ? $signed(_GEN_451) : $signed(_GEN_435); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_468 = activeSums_10 ? $signed(_GEN_452) : $signed(_GEN_436); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_469 = activeSums_10 ? $signed(_GEN_453) : $signed(_GEN_437); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_470 = activeSums_10 ? $signed(_GEN_454) : $signed(_GEN_438); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_471 = activeSums_10 ? $signed(_GEN_455) : $signed(_GEN_439); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_472 = activeSums_10 ? $signed(_GEN_456) : $signed(_GEN_440); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_473 = activeSums_10 ? $signed(_GEN_457) : $signed(_GEN_441); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_474 = activeSums_10 ? $signed(_GEN_458) : $signed(_GEN_442); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_475 = activeSums_10 ? $signed(_GEN_459) : $signed(_GEN_443); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_476 = activeSums_10 ? $signed(_GEN_460) : $signed(_GEN_444); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_477 = activeSums_10 ? $signed(_GEN_461) : $signed(_GEN_445); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_478 = activeSums_10 ? $signed(_GEN_462) : $signed(_GEN_446); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_11 = _T_588; // @[CFARCoreWithASR.scala 110:29]
  assign _T_886 = 4'hb >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_479 = 4'h0 == _T_886 ? $signed(max_11) : $signed(_GEN_463); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_480 = 4'h1 == _T_886 ? $signed(max_11) : $signed(_GEN_464); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_481 = 4'h2 == _T_886 ? $signed(max_11) : $signed(_GEN_465); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_482 = 4'h3 == _T_886 ? $signed(max_11) : $signed(_GEN_466); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_483 = 4'h4 == _T_886 ? $signed(max_11) : $signed(_GEN_467); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_484 = 4'h5 == _T_886 ? $signed(max_11) : $signed(_GEN_468); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_485 = 4'h6 == _T_886 ? $signed(max_11) : $signed(_GEN_469); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_486 = 4'h7 == _T_886 ? $signed(max_11) : $signed(_GEN_470); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_487 = 4'h8 == _T_886 ? $signed(max_11) : $signed(_GEN_471); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_488 = 4'h9 == _T_886 ? $signed(max_11) : $signed(_GEN_472); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_489 = 4'ha == _T_886 ? $signed(max_11) : $signed(_GEN_473); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_490 = 4'hb == _T_886 ? $signed(max_11) : $signed(_GEN_474); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_491 = 4'hc == _T_886 ? $signed(max_11) : $signed(_GEN_475); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_492 = 4'hd == _T_886 ? $signed(max_11) : $signed(_GEN_476); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_493 = 4'he == _T_886 ? $signed(max_11) : $signed(_GEN_477); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_494 = 4'hf == _T_886 ? $signed(max_11) : $signed(_GEN_478); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_495 = activeSums_11 ? $signed(_GEN_479) : $signed(_GEN_463); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_496 = activeSums_11 ? $signed(_GEN_480) : $signed(_GEN_464); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_497 = activeSums_11 ? $signed(_GEN_481) : $signed(_GEN_465); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_498 = activeSums_11 ? $signed(_GEN_482) : $signed(_GEN_466); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_499 = activeSums_11 ? $signed(_GEN_483) : $signed(_GEN_467); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_500 = activeSums_11 ? $signed(_GEN_484) : $signed(_GEN_468); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_501 = activeSums_11 ? $signed(_GEN_485) : $signed(_GEN_469); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_502 = activeSums_11 ? $signed(_GEN_486) : $signed(_GEN_470); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_503 = activeSums_11 ? $signed(_GEN_487) : $signed(_GEN_471); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_504 = activeSums_11 ? $signed(_GEN_488) : $signed(_GEN_472); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_505 = activeSums_11 ? $signed(_GEN_489) : $signed(_GEN_473); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_506 = activeSums_11 ? $signed(_GEN_490) : $signed(_GEN_474); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_507 = activeSums_11 ? $signed(_GEN_491) : $signed(_GEN_475); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_508 = activeSums_11 ? $signed(_GEN_492) : $signed(_GEN_476); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_509 = activeSums_11 ? $signed(_GEN_493) : $signed(_GEN_477); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_510 = activeSums_11 ? $signed(_GEN_494) : $signed(_GEN_478); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_12 = _T_633; // @[CFARCoreWithASR.scala 110:29]
  assign _T_888 = 4'hc >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_511 = 4'h0 == _T_888 ? $signed(max_12) : $signed(_GEN_495); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_512 = 4'h1 == _T_888 ? $signed(max_12) : $signed(_GEN_496); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_513 = 4'h2 == _T_888 ? $signed(max_12) : $signed(_GEN_497); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_514 = 4'h3 == _T_888 ? $signed(max_12) : $signed(_GEN_498); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_515 = 4'h4 == _T_888 ? $signed(max_12) : $signed(_GEN_499); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_516 = 4'h5 == _T_888 ? $signed(max_12) : $signed(_GEN_500); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_517 = 4'h6 == _T_888 ? $signed(max_12) : $signed(_GEN_501); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_518 = 4'h7 == _T_888 ? $signed(max_12) : $signed(_GEN_502); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_519 = 4'h8 == _T_888 ? $signed(max_12) : $signed(_GEN_503); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_520 = 4'h9 == _T_888 ? $signed(max_12) : $signed(_GEN_504); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_521 = 4'ha == _T_888 ? $signed(max_12) : $signed(_GEN_505); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_522 = 4'hb == _T_888 ? $signed(max_12) : $signed(_GEN_506); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_523 = 4'hc == _T_888 ? $signed(max_12) : $signed(_GEN_507); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_524 = 4'hd == _T_888 ? $signed(max_12) : $signed(_GEN_508); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_525 = 4'he == _T_888 ? $signed(max_12) : $signed(_GEN_509); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_526 = 4'hf == _T_888 ? $signed(max_12) : $signed(_GEN_510); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_527 = activeSums_12 ? $signed(_GEN_511) : $signed(_GEN_495); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_528 = activeSums_12 ? $signed(_GEN_512) : $signed(_GEN_496); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_529 = activeSums_12 ? $signed(_GEN_513) : $signed(_GEN_497); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_530 = activeSums_12 ? $signed(_GEN_514) : $signed(_GEN_498); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_531 = activeSums_12 ? $signed(_GEN_515) : $signed(_GEN_499); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_532 = activeSums_12 ? $signed(_GEN_516) : $signed(_GEN_500); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_533 = activeSums_12 ? $signed(_GEN_517) : $signed(_GEN_501); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_534 = activeSums_12 ? $signed(_GEN_518) : $signed(_GEN_502); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_535 = activeSums_12 ? $signed(_GEN_519) : $signed(_GEN_503); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_536 = activeSums_12 ? $signed(_GEN_520) : $signed(_GEN_504); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_537 = activeSums_12 ? $signed(_GEN_521) : $signed(_GEN_505); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_538 = activeSums_12 ? $signed(_GEN_522) : $signed(_GEN_506); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_539 = activeSums_12 ? $signed(_GEN_523) : $signed(_GEN_507); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_540 = activeSums_12 ? $signed(_GEN_524) : $signed(_GEN_508); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_541 = activeSums_12 ? $signed(_GEN_525) : $signed(_GEN_509); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_542 = activeSums_12 ? $signed(_GEN_526) : $signed(_GEN_510); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_13 = _T_678; // @[CFARCoreWithASR.scala 110:29]
  assign _T_890 = 4'hd >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_543 = 4'h0 == _T_890 ? $signed(max_13) : $signed(_GEN_527); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_544 = 4'h1 == _T_890 ? $signed(max_13) : $signed(_GEN_528); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_545 = 4'h2 == _T_890 ? $signed(max_13) : $signed(_GEN_529); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_546 = 4'h3 == _T_890 ? $signed(max_13) : $signed(_GEN_530); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_547 = 4'h4 == _T_890 ? $signed(max_13) : $signed(_GEN_531); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_548 = 4'h5 == _T_890 ? $signed(max_13) : $signed(_GEN_532); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_549 = 4'h6 == _T_890 ? $signed(max_13) : $signed(_GEN_533); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_550 = 4'h7 == _T_890 ? $signed(max_13) : $signed(_GEN_534); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_551 = 4'h8 == _T_890 ? $signed(max_13) : $signed(_GEN_535); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_552 = 4'h9 == _T_890 ? $signed(max_13) : $signed(_GEN_536); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_553 = 4'ha == _T_890 ? $signed(max_13) : $signed(_GEN_537); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_554 = 4'hb == _T_890 ? $signed(max_13) : $signed(_GEN_538); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_555 = 4'hc == _T_890 ? $signed(max_13) : $signed(_GEN_539); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_556 = 4'hd == _T_890 ? $signed(max_13) : $signed(_GEN_540); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_557 = 4'he == _T_890 ? $signed(max_13) : $signed(_GEN_541); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_558 = 4'hf == _T_890 ? $signed(max_13) : $signed(_GEN_542); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_559 = activeSums_13 ? $signed(_GEN_543) : $signed(_GEN_527); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_560 = activeSums_13 ? $signed(_GEN_544) : $signed(_GEN_528); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_561 = activeSums_13 ? $signed(_GEN_545) : $signed(_GEN_529); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_562 = activeSums_13 ? $signed(_GEN_546) : $signed(_GEN_530); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_563 = activeSums_13 ? $signed(_GEN_547) : $signed(_GEN_531); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_564 = activeSums_13 ? $signed(_GEN_548) : $signed(_GEN_532); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_565 = activeSums_13 ? $signed(_GEN_549) : $signed(_GEN_533); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_566 = activeSums_13 ? $signed(_GEN_550) : $signed(_GEN_534); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_567 = activeSums_13 ? $signed(_GEN_551) : $signed(_GEN_535); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_568 = activeSums_13 ? $signed(_GEN_552) : $signed(_GEN_536); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_569 = activeSums_13 ? $signed(_GEN_553) : $signed(_GEN_537); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_570 = activeSums_13 ? $signed(_GEN_554) : $signed(_GEN_538); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_571 = activeSums_13 ? $signed(_GEN_555) : $signed(_GEN_539); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_572 = activeSums_13 ? $signed(_GEN_556) : $signed(_GEN_540); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_573 = activeSums_13 ? $signed(_GEN_557) : $signed(_GEN_541); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_574 = activeSums_13 ? $signed(_GEN_558) : $signed(_GEN_542); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_14 = _T_721; // @[CFARCoreWithASR.scala 110:29]
  assign _T_892 = 4'he >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_575 = 4'h0 == _T_892 ? $signed(max_14) : $signed(_GEN_559); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_576 = 4'h1 == _T_892 ? $signed(max_14) : $signed(_GEN_560); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_577 = 4'h2 == _T_892 ? $signed(max_14) : $signed(_GEN_561); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_578 = 4'h3 == _T_892 ? $signed(max_14) : $signed(_GEN_562); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_579 = 4'h4 == _T_892 ? $signed(max_14) : $signed(_GEN_563); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_580 = 4'h5 == _T_892 ? $signed(max_14) : $signed(_GEN_564); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_581 = 4'h6 == _T_892 ? $signed(max_14) : $signed(_GEN_565); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_582 = 4'h7 == _T_892 ? $signed(max_14) : $signed(_GEN_566); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_583 = 4'h8 == _T_892 ? $signed(max_14) : $signed(_GEN_567); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_584 = 4'h9 == _T_892 ? $signed(max_14) : $signed(_GEN_568); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_585 = 4'ha == _T_892 ? $signed(max_14) : $signed(_GEN_569); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_586 = 4'hb == _T_892 ? $signed(max_14) : $signed(_GEN_570); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_587 = 4'hc == _T_892 ? $signed(max_14) : $signed(_GEN_571); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_588 = 4'hd == _T_892 ? $signed(max_14) : $signed(_GEN_572); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_589 = 4'he == _T_892 ? $signed(max_14) : $signed(_GEN_573); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_590 = 4'hf == _T_892 ? $signed(max_14) : $signed(_GEN_574); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_591 = activeSums_14 ? $signed(_GEN_575) : $signed(_GEN_559); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_592 = activeSums_14 ? $signed(_GEN_576) : $signed(_GEN_560); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_593 = activeSums_14 ? $signed(_GEN_577) : $signed(_GEN_561); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_594 = activeSums_14 ? $signed(_GEN_578) : $signed(_GEN_562); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_595 = activeSums_14 ? $signed(_GEN_579) : $signed(_GEN_563); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_596 = activeSums_14 ? $signed(_GEN_580) : $signed(_GEN_564); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_597 = activeSums_14 ? $signed(_GEN_581) : $signed(_GEN_565); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_598 = activeSums_14 ? $signed(_GEN_582) : $signed(_GEN_566); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_599 = activeSums_14 ? $signed(_GEN_583) : $signed(_GEN_567); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_600 = activeSums_14 ? $signed(_GEN_584) : $signed(_GEN_568); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_601 = activeSums_14 ? $signed(_GEN_585) : $signed(_GEN_569); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_602 = activeSums_14 ? $signed(_GEN_586) : $signed(_GEN_570); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_603 = activeSums_14 ? $signed(_GEN_587) : $signed(_GEN_571); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_604 = activeSums_14 ? $signed(_GEN_588) : $signed(_GEN_572); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_605 = activeSums_14 ? $signed(_GEN_589) : $signed(_GEN_573); // @[CFARCoreWithASR.scala 200:32]
  assign _GEN_606 = activeSums_14 ? $signed(_GEN_590) : $signed(_GEN_574); // @[CFARCoreWithASR.scala 200:32]
  assign activeSums_15 = _T_764; // @[CFARCoreWithASR.scala 110:29]
  assign _T_894 = 4'hf >> diffInSubSize; // @[CFARCoreWithASR.scala 201:29]
  assign _GEN_607 = 4'h0 == _T_894 ? $signed(max_15) : $signed(_GEN_591); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_608 = 4'h1 == _T_894 ? $signed(max_15) : $signed(_GEN_592); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_609 = 4'h2 == _T_894 ? $signed(max_15) : $signed(_GEN_593); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_610 = 4'h3 == _T_894 ? $signed(max_15) : $signed(_GEN_594); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_611 = 4'h4 == _T_894 ? $signed(max_15) : $signed(_GEN_595); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_612 = 4'h5 == _T_894 ? $signed(max_15) : $signed(_GEN_596); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_613 = 4'h6 == _T_894 ? $signed(max_15) : $signed(_GEN_597); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_614 = 4'h7 == _T_894 ? $signed(max_15) : $signed(_GEN_598); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_615 = 4'h8 == _T_894 ? $signed(max_15) : $signed(_GEN_599); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_616 = 4'h9 == _T_894 ? $signed(max_15) : $signed(_GEN_600); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_617 = 4'ha == _T_894 ? $signed(max_15) : $signed(_GEN_601); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_618 = 4'hb == _T_894 ? $signed(max_15) : $signed(_GEN_602); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_619 = 4'hc == _T_894 ? $signed(max_15) : $signed(_GEN_603); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_620 = 4'hd == _T_894 ? $signed(max_15) : $signed(_GEN_604); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_621 = 4'he == _T_894 ? $signed(max_15) : $signed(_GEN_605); // @[CFARCoreWithASR.scala 202:27]
  assign _GEN_622 = 4'hf == _T_894 ? $signed(max_15) : $signed(_GEN_606); // @[CFARCoreWithASR.scala 202:27]
  assign _T_908 = io_windowCells >> _T_811; // @[CFARCoreWithASR.scala 209:46]
  assign clutterRepr = $signed(minCircuit_io_out) >>> _T_811; // @[FixedPointTypeClass.scala 118:51]
  assign _T_924 = cntIn + 9'h1; // @[CFARCoreWithASR.scala 216:20]
  assign _T_926 = latency - 9'h1; // @[CFARCoreWithASR.scala 218:28]
  assign _T_927 = cntIn == _T_926; // @[CFARCoreWithASR.scala 218:15]
  assign _T_929 = _T_927 & _T_114; // @[CFARCoreWithASR.scala 218:35]
  assign _GEN_640 = _T_929 | initialInDone; // @[CFARCoreWithASR.scala 218:52]
  assign _T_930 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_931 = io_lastOut & _T_930; // @[CFARCoreWithASR.scala 222:20]
  assign _T_934 = cntOut + 9'h1; // @[CFARCoreWithASR.scala 226:22]
  assign _T_936 = io_fftWin - 10'h1; // @[CFARCoreWithASR.scala 228:31]
  assign _GEN_916 = {{1'd0}, cntOut}; // @[CFARCoreWithASR.scala 228:16]
  assign _T_937 = _GEN_916 == _T_936; // @[CFARCoreWithASR.scala 228:16]
  assign _T_939 = _T_937 & _T_930; // @[CFARCoreWithASR.scala 228:38]
  assign _T_942 = _T_939 | _T_931; // @[CFARCoreWithASR.scala 228:55]
  assign _GEN_644 = io_lastIn | flushing; // @[CFARCoreWithASR.scala 232:20]
  assign leftThr = $signed(sumSubLaggs_0) >>> io_divSum; // @[FixedPointTypeClass.scala 118:51]
  assign rightThr = $signed(sumSubLeads_0) >>> io_divSum; // @[FixedPointTypeClass.scala 118:51]
  assign _T_944 = $signed(leftThr) > $signed(rightThr); // @[FixedPointTypeClass.scala 55:59]
  assign greatestOf = _T_944 ? $signed(leftThr) : $signed(rightThr); // @[CFARCoreWithASR.scala 289:23]
  assign _T_945 = $signed(leftThr) < $signed(rightThr); // @[FixedPointTypeClass.scala 53:59]
  assign smallestOf = _T_945 ? $signed(leftThr) : $signed(rightThr); // @[CFARCoreWithASR.scala 290:23]
  assign _T_948 = $signed(rightThr) + $signed(leftThr); // @[FixedPointTypeClass.scala 20:58]
  assign _T_949 = _T_948[19:1]; // @[FixedPointTypeClass.scala 117:50]
  assign _T_950 = 2'h3 == io_cfarMode; // @[Mux.scala 68:19]
  assign _T_951 = _T_950 ? $signed(clutterRepr) : $signed(smallestOf); // @[Mux.scala 68:16]
  assign _T_952 = 2'h2 == io_cfarMode; // @[Mux.scala 68:19]
  assign _T_953 = _T_952 ? $signed(smallestOf) : $signed(_T_951); // @[Mux.scala 68:16]
  assign _T_954 = 2'h1 == io_cfarMode; // @[Mux.scala 68:19]
  assign _T_955 = _T_954 ? $signed(greatestOf) : $signed(_T_953); // @[Mux.scala 68:16]
  assign _T_956 = 2'h0 == io_cfarMode; // @[Mux.scala 68:19]
  assign thrByModes = _T_956 ? $signed({{1{_T_949[18]}},_T_949}) : $signed(_T_955); // @[Mux.scala 68:16]
  assign _T_957 = ~laggWindow_io_regFull; // @[CFARCoreWithASR.scala 300:9]
  assign _T_958 = laggWindow_io_out_ready & laggWindow_io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_959 = _T_957 & _T_958; // @[CFARCoreWithASR.scala 300:34]
  assign _GEN_651 = _T_959 | enableRightThr; // @[CFARCoreWithASR.scala 300:63]
  assign _T_960 = laggWindow_io_regFull & leadWindow_io_regFull; // @[CFARCoreWithASR.scala 313:50]
  assign _T_961 = ~leadWindow_io_regFull; // @[CFARCoreWithASR.scala 315:60]
  assign _T_962 = enableRightThr | _T_961; // @[CFARCoreWithASR.scala 315:57]
  assign _T_963 = enableRightThr ? $signed(rightThr) : $signed(leftThr); // @[CFARCoreWithASR.scala 315:87]
  assign _T_964 = _T_962 ? $signed(_T_963) : $signed(thrByModes); // @[CFARCoreWithASR.scala 315:41]
  assign thrWithoutScaling = _T_960 ? $signed(thrByModes) : $signed(_T_964); // @[CFARCoreWithASR.scala 313:27]
  assign _GEN_917 = {{4{io_thresholdScaler[15]}},io_thresholdScaler}; // @[FixedPointTypeClass.scala 211:35]
  assign threshold = _T_966[35:13]; // @[FixedPointTypeClass.scala 153:43]
  assign _T_967 = io_guardCells == 4'h0; // @[CFARCoreWithASR.scala 394:53]
  assign _T_969 = io_windowCells - 7'h1; // @[CFARCoreWithASR.scala 394:103]
  assign _T_972 = io_guardCells - 4'h1; // @[CFARCoreWithASR.scala 394:150]
  assign _GEN_655 = laggWindow_io_parallelOut_0; // @[CFARCoreWithASR.scala 394:38]
  assign _GEN_719 = laggGuard_io_parallelOut_0; // @[CFARCoreWithASR.scala 394:38]
  assign _T_977 = $signed(cutDelayed) > $signed(leftNeighb); // @[FixedPointTypeClass.scala 55:59]
  assign _T_978 = $signed(cutDelayed) > $signed(rightNeighb); // @[FixedPointTypeClass.scala 55:59]
  assign isLocalMax = _T_977 & _T_978; // @[CFARCoreWithASR.scala 396:44]
  assign _GEN_918 = {$signed(cutDelayed), 1'h0}; // @[FixedPointTypeClass.scala 55:59]
  assign _GEN_919 = {{6{_GEN_918[16]}},_GEN_918}; // @[FixedPointTypeClass.scala 55:59]
  assign isPeak = $signed(_GEN_919) > $signed(threshold); // @[FixedPointTypeClass.scala 55:59]
  assign _T_979 = ~initialInDone; // @[CFARCoreWithASR.scala 418:20]
  assign _T_980 = ~flushingDelayed; // @[CFARCoreWithASR.scala 418:54]
  assign _T_981 = io_out_ready & _T_980; // @[CFARCoreWithASR.scala 418:51]
  assign _T_987 = flushingDelayed & _T_986; // @[CFARCoreWithASR.scala 419:121]
  assign _T_989 = isPeak & isLocalMax; // @[CFARCoreWithASR.scala 430:65]
  assign _T_995 = flushingDelayed & _T_994; // @[CFARCoreWithASR.scala 435:121]
  assign io_in_ready = _T_979 | _T_981; // @[CFARCoreWithASR.scala 44:20 CFARCoreWithASR.scala 418:17]
  assign io_out_valid = Queue_io_deq_valid; // @[CFARCoreWithASR.scala 446:18]
  assign io_out_bits_peak = Queue_io_deq_bits_peak; // @[CFARCoreWithASR.scala 443:22]
  assign io_out_bits_cut = Queue_io_deq_bits_cut; // @[CFARCoreWithASR.scala 442:27]
  assign io_out_bits_threshold = Queue_io_deq_bits_threshold; // @[CFARCoreWithASR.scala 444:27]
  assign io_lastOut = Queue_1_io_deq_bits; // @[CFARCoreWithASR.scala 439:16]
  assign io_fftBin = cntOut; // @[CFARCoreWithASR.scala 447:15]
  assign laggWindow_clock = clock;
  assign laggWindow_reset = reset;
  assign laggWindow_io_depth = io_windowCells; // @[CFARCoreWithASR.scala 45:23]
  assign laggWindow_io_in_valid = io_in_valid; // @[CFARCoreWithASR.scala 44:20]
  assign laggWindow_io_in_bits = io_in_bits; // @[CFARCoreWithASR.scala 44:20]
  assign laggWindow_io_lastIn = io_lastIn; // @[CFARCoreWithASR.scala 46:24]
  assign laggWindow_io_out_ready = laggGuard_io_in_ready; // @[CFARCoreWithASR.scala 59:19]
  assign laggGuard_clock = clock;
  assign laggGuard_reset = reset;
  assign laggGuard_io_depth = io_guardCells; // @[CFARCoreWithASR.scala 61:23]
  assign laggGuard_io_in_valid = laggWindow_io_out_valid; // @[CFARCoreWithASR.scala 59:19]
  assign laggGuard_io_in_bits = laggWindow_io_out_bits; // @[CFARCoreWithASR.scala 59:19]
  assign laggGuard_io_lastIn = laggWindow_io_lastOut; // @[CFARCoreWithASR.scala 60:23]
  assign laggGuard_io_out_ready = cellUnderTest_io_in_ready; // @[CFARCoreWithASR.scala 64:23]
  assign cellUnderTest_clock = clock;
  assign cellUnderTest_reset = reset;
  assign cellUnderTest_io_in_valid = laggGuard_io_out_valid; // @[CFARCoreWithASR.scala 64:23]
  assign cellUnderTest_io_in_bits = laggGuard_io_out_bits; // @[CFARCoreWithASR.scala 64:23]
  assign cellUnderTest_io_lastIn = laggGuard_io_lastOut; // @[CFARCoreWithASR.scala 65:27]
  assign cellUnderTest_io_out_ready = leadWindow_io_regFull ? leadWindow_io_in_ready : io_out_ready; // @[CFARCoreWithASR.scala 69:19 CFARCoreWithASR.scala 83:30]
  assign leadGuard_clock = clock;
  assign leadGuard_reset = reset;
  assign leadGuard_io_depth = io_guardCells; // @[CFARCoreWithASR.scala 70:22]
  assign leadGuard_io_in_valid = cellUnderTest_io_out_valid; // @[CFARCoreWithASR.scala 69:19]
  assign leadGuard_io_in_bits = cellUnderTest_io_out_bits; // @[CFARCoreWithASR.scala 69:19]
  assign leadGuard_io_lastIn = cellUnderTest_io_lastOut; // @[CFARCoreWithASR.scala 71:23]
  assign leadGuard_io_out_ready = leadWindow_io_in_ready; // @[CFARCoreWithASR.scala 72:26 CFARCoreWithASR.scala 76:20]
  assign leadWindow_clock = clock;
  assign leadWindow_reset = reset;
  assign leadWindow_io_depth = io_windowCells; // @[CFARCoreWithASR.scala 75:23]
  assign leadWindow_io_in_valid = leadGuard_io_out_valid; // @[CFARCoreWithASR.scala 76:20]
  assign leadWindow_io_in_bits = leadGuard_io_out_bits; // @[CFARCoreWithASR.scala 76:20]
  assign leadWindow_io_lastIn = leadGuard_io_lastOut; // @[CFARCoreWithASR.scala 84:24]
  assign leadWindow_io_out_ready = io_out_ready; // @[CFARCoreWithASR.scala 79:27]
  assign minCircuit_clock = clock;
  assign minCircuit_io_in_0 = activeSums_15 ? $signed(_GEN_607) : $signed(_GEN_591); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_1 = activeSums_15 ? $signed(_GEN_608) : $signed(_GEN_592); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_2 = activeSums_15 ? $signed(_GEN_609) : $signed(_GEN_593); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_3 = activeSums_15 ? $signed(_GEN_610) : $signed(_GEN_594); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_4 = activeSums_15 ? $signed(_GEN_611) : $signed(_GEN_595); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_5 = activeSums_15 ? $signed(_GEN_612) : $signed(_GEN_596); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_6 = activeSums_15 ? $signed(_GEN_613) : $signed(_GEN_597); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_7 = activeSums_15 ? $signed(_GEN_614) : $signed(_GEN_598); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_8 = activeSums_15 ? $signed(_GEN_615) : $signed(_GEN_599); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_9 = activeSums_15 ? $signed(_GEN_616) : $signed(_GEN_600); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_10 = activeSums_15 ? $signed(_GEN_617) : $signed(_GEN_601); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_11 = activeSums_15 ? $signed(_GEN_618) : $signed(_GEN_602); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_12 = activeSums_15 ? $signed(_GEN_619) : $signed(_GEN_603); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_13 = activeSums_15 ? $signed(_GEN_620) : $signed(_GEN_604); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_14 = activeSums_15 ? $signed(_GEN_621) : $signed(_GEN_605); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_in_15 = activeSums_15 ? $signed(_GEN_622) : $signed(_GEN_606); // @[CFARCoreWithASR.scala 208:20]
  assign minCircuit_io_inSize = _T_908[4:0]; // @[CFARCoreWithASR.scala 209:28]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_985 | _T_987; // @[CFARCoreWithASR.scala 419:28]
  assign Queue_io_enq_bits_peak = io_peakGrouping ? _T_989 : isPeak; // @[CFARCoreWithASR.scala 430:34]
  assign Queue_io_enq_bits_cut = cutDelayed; // @[CFARCoreWithASR.scala 422:37]
  assign _GEN_921 = threshold[22:1]; // @[CFARCoreWithASR.scala 423:37]
  assign Queue_io_enq_bits_threshold = _GEN_921[15:0]; // @[CFARCoreWithASR.scala 423:37]
  assign Queue_io_deq_ready = io_out_ready; // @[CFARCoreWithASR.scala 432:28]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_993 | _T_995; // @[CFARCoreWithASR.scala 435:28]
  assign Queue_1_io_enq_bits = lastOut; // @[CFARCoreWithASR.scala 436:27]
  assign Queue_1_io_deq_ready = io_out_ready; // @[CFARCoreWithASR.scala 438:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flushing = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntIn = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cntOut = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  initialInDone = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  lastOut = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sumSubLaggs_0 = _RAND_5[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sumSubLaggs_1 = _RAND_6[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sumSubLaggs_2 = _RAND_7[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sumSubLaggs_3 = _RAND_8[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sumSubLaggs_4 = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  sumSubLaggs_5 = _RAND_10[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  sumSubLaggs_6 = _RAND_11[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  sumSubLaggs_7 = _RAND_12[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  sumSubLaggs_8 = _RAND_13[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sumSubLaggs_9 = _RAND_14[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sumSubLaggs_10 = _RAND_15[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sumSubLaggs_11 = _RAND_16[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sumSubLaggs_12 = _RAND_17[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sumSubLaggs_13 = _RAND_18[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  sumSubLaggs_14 = _RAND_19[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  sumSubLaggs_15 = _RAND_20[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  sumSubLeads_0 = _RAND_21[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  sumSubLeads_1 = _RAND_22[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sumSubLeads_2 = _RAND_23[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sumSubLeads_3 = _RAND_24[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sumSubLeads_4 = _RAND_25[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sumSubLeads_5 = _RAND_26[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sumSubLeads_6 = _RAND_27[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  sumSubLeads_7 = _RAND_28[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  sumSubLeads_8 = _RAND_29[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  sumSubLeads_9 = _RAND_30[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  sumSubLeads_10 = _RAND_31[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sumSubLeads_11 = _RAND_32[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sumSubLeads_12 = _RAND_33[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sumSubLeads_13 = _RAND_34[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sumSubLeads_14 = _RAND_35[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sumSubLeads_15 = _RAND_36[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  flushingDelayed = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  enableRightThr = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_966 = _RAND_39[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  cutDelayed = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  leftNeighb = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  rightNeighb = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_985 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_986 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_993 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_994 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flushing <= 1'h0;
    end else if (lastOut) begin
      flushing <= 1'h0;
    end else begin
      flushing <= _GEN_644;
    end
    if (reset) begin
      cntIn <= 9'h0;
    end else if (_T_931) begin
      cntIn <= 9'h0;
    end else if (_T_114) begin
      cntIn <= _T_924;
    end
    if (reset) begin
      cntOut <= 9'h0;
    end else if (_T_942) begin
      cntOut <= 9'h0;
    end else if (_T_930) begin
      cntOut <= _T_934;
    end
    if (reset) begin
      initialInDone <= 1'h0;
    end else if (lastOut) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_640;
    end
    lastOut <= cellUnderTest_io_lastOut;
    if (reset) begin
      sumSubLaggs_0 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_0 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_115) begin
        sumSubLaggs_0 <= _T_121;
      end else begin
        sumSubLaggs_0 <= _T_118;
      end
    end
    if (reset) begin
      sumSubLaggs_1 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_1 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_156) begin
        sumSubLaggs_1 <= _T_162;
      end else if (maybeFullLagg_0) begin
        sumSubLaggs_1 <= _T_159;
      end
    end
    if (reset) begin
      sumSubLaggs_2 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_2 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_201) begin
        sumSubLaggs_2 <= _T_207;
      end else if (maybeFullLagg_1) begin
        sumSubLaggs_2 <= _T_204;
      end
    end
    if (reset) begin
      sumSubLaggs_3 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_3 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_242) begin
        sumSubLaggs_3 <= _T_248;
      end else if (maybeFullLagg_2) begin
        sumSubLaggs_3 <= _T_245;
      end
    end
    if (reset) begin
      sumSubLaggs_4 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_4 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_291) begin
        sumSubLaggs_4 <= _T_297;
      end else if (maybeFullLagg_3) begin
        sumSubLaggs_4 <= _T_294;
      end
    end
    if (reset) begin
      sumSubLaggs_5 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_5 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_332) begin
        sumSubLaggs_5 <= _T_338;
      end else if (maybeFullLagg_4) begin
        sumSubLaggs_5 <= _T_335;
      end
    end
    if (reset) begin
      sumSubLaggs_6 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_6 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_377) begin
        sumSubLaggs_6 <= _T_383;
      end else if (maybeFullLagg_5) begin
        sumSubLaggs_6 <= _T_380;
      end
    end
    if (reset) begin
      sumSubLaggs_7 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_7 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_418) begin
        sumSubLaggs_7 <= _T_424;
      end else if (maybeFullLagg_6) begin
        sumSubLaggs_7 <= _T_421;
      end
    end
    if (reset) begin
      sumSubLaggs_8 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_8 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_471) begin
        sumSubLaggs_8 <= _T_477;
      end else if (maybeFullLagg_7) begin
        sumSubLaggs_8 <= _T_474;
      end
    end
    if (reset) begin
      sumSubLaggs_9 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_9 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_512) begin
        sumSubLaggs_9 <= _T_518;
      end else if (maybeFullLagg_8) begin
        sumSubLaggs_9 <= _T_515;
      end
    end
    if (reset) begin
      sumSubLaggs_10 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_10 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_557) begin
        sumSubLaggs_10 <= _T_563;
      end else if (maybeFullLagg_9) begin
        sumSubLaggs_10 <= _T_560;
      end
    end
    if (reset) begin
      sumSubLaggs_11 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_11 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_598) begin
        sumSubLaggs_11 <= _T_604;
      end else if (maybeFullLagg_10) begin
        sumSubLaggs_11 <= _T_601;
      end
    end
    if (reset) begin
      sumSubLaggs_12 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_12 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_647) begin
        sumSubLaggs_12 <= _T_653;
      end else if (maybeFullLagg_11) begin
        sumSubLaggs_12 <= _T_650;
      end
    end
    if (reset) begin
      sumSubLaggs_13 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_13 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_688) begin
        sumSubLaggs_13 <= _T_694;
      end else if (maybeFullLagg_12) begin
        sumSubLaggs_13 <= _T_691;
      end
    end
    if (reset) begin
      sumSubLaggs_14 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_14 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_733) begin
        sumSubLaggs_14 <= _T_739;
      end else if (maybeFullLagg_13) begin
        sumSubLaggs_14 <= _T_736;
      end
    end
    if (reset) begin
      sumSubLaggs_15 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLaggs_15 <= 20'sh0;
    end else if (_T_114) begin
      if (_T_774) begin
        sumSubLaggs_15 <= _T_780;
      end else if (maybeFullLagg_14) begin
        sumSubLaggs_15 <= _T_777;
      end
    end
    if (reset) begin
      sumSubLeads_0 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_0 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_130) begin
        sumSubLeads_0 <= _T_136;
      end else begin
        sumSubLeads_0 <= _T_133;
      end
    end
    if (reset) begin
      sumSubLeads_1 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_1 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_171) begin
        sumSubLeads_1 <= _T_177;
      end else if (maybeFullLead_0) begin
        sumSubLeads_1 <= _T_174;
      end
    end
    if (reset) begin
      sumSubLeads_2 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_2 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_216) begin
        sumSubLeads_2 <= _T_222;
      end else if (maybeFullLead_1) begin
        sumSubLeads_2 <= _T_219;
      end
    end
    if (reset) begin
      sumSubLeads_3 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_3 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_257) begin
        sumSubLeads_3 <= _T_263;
      end else if (maybeFullLead_2) begin
        sumSubLeads_3 <= _T_260;
      end
    end
    if (reset) begin
      sumSubLeads_4 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_4 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_306) begin
        sumSubLeads_4 <= _T_312;
      end else if (maybeFullLead_3) begin
        sumSubLeads_4 <= _T_309;
      end
    end
    if (reset) begin
      sumSubLeads_5 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_5 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_347) begin
        sumSubLeads_5 <= _T_353;
      end else if (maybeFullLead_4) begin
        sumSubLeads_5 <= _T_350;
      end
    end
    if (reset) begin
      sumSubLeads_6 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_6 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_392) begin
        sumSubLeads_6 <= _T_398;
      end else if (maybeFullLead_5) begin
        sumSubLeads_6 <= _T_395;
      end
    end
    if (reset) begin
      sumSubLeads_7 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_7 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_433) begin
        sumSubLeads_7 <= _T_439;
      end else if (maybeFullLead_6) begin
        sumSubLeads_7 <= _T_436;
      end
    end
    if (reset) begin
      sumSubLeads_8 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_8 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_486) begin
        sumSubLeads_8 <= _T_492;
      end else if (maybeFullLead_7) begin
        sumSubLeads_8 <= _T_489;
      end
    end
    if (reset) begin
      sumSubLeads_9 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_9 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_527) begin
        sumSubLeads_9 <= _T_533;
      end else if (maybeFullLead_8) begin
        sumSubLeads_9 <= _T_530;
      end
    end
    if (reset) begin
      sumSubLeads_10 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_10 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_572) begin
        sumSubLeads_10 <= _T_578;
      end else if (maybeFullLead_9) begin
        sumSubLeads_10 <= _T_575;
      end
    end
    if (reset) begin
      sumSubLeads_11 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_11 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_613) begin
        sumSubLeads_11 <= _T_619;
      end else if (maybeFullLead_10) begin
        sumSubLeads_11 <= _T_616;
      end
    end
    if (reset) begin
      sumSubLeads_12 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_12 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_662) begin
        sumSubLeads_12 <= _T_668;
      end else if (maybeFullLead_11) begin
        sumSubLeads_12 <= _T_665;
      end
    end
    if (reset) begin
      sumSubLeads_13 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_13 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_703) begin
        sumSubLeads_13 <= _T_709;
      end else if (maybeFullLead_12) begin
        sumSubLeads_13 <= _T_706;
      end
    end
    if (reset) begin
      sumSubLeads_14 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_14 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_748) begin
        sumSubLeads_14 <= _T_754;
      end else if (maybeFullLead_13) begin
        sumSubLeads_14 <= _T_751;
      end
    end
    if (reset) begin
      sumSubLeads_15 <= 20'sh0;
    end else if (io_lastOut) begin
      sumSubLeads_15 <= 20'sh0;
    end else if (_T_129) begin
      if (_T_789) begin
        sumSubLeads_15 <= _T_795;
      end else if (maybeFullLead_14) begin
        sumSubLeads_15 <= _T_792;
      end
    end
    if (reset) begin
      flushingDelayed <= 1'h0;
    end else if (io_lastOut) begin
      flushingDelayed <= 1'h0;
    end else begin
      flushingDelayed <= flushing;
    end
    if (reset) begin
      enableRightThr <= 1'h0;
    end else if (io_lastOut) begin
      enableRightThr <= 1'h0;
    end else begin
      enableRightThr <= _GEN_651;
    end
    _T_966 <= $signed(thrWithoutScaling) * $signed(_GEN_917);
    cutDelayed <= cellUnderTest_io_out_bits;
    if (_T_967) begin
      if (6'h3f == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_63;
      end else if (6'h3e == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_62;
      end else if (6'h3d == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_61;
      end else if (6'h3c == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_60;
      end else if (6'h3b == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_59;
      end else if (6'h3a == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_58;
      end else if (6'h39 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_57;
      end else if (6'h38 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_56;
      end else if (6'h37 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_55;
      end else if (6'h36 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_54;
      end else if (6'h35 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_53;
      end else if (6'h34 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_52;
      end else if (6'h33 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_51;
      end else if (6'h32 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_50;
      end else if (6'h31 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_49;
      end else if (6'h30 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_48;
      end else if (6'h2f == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_47;
      end else if (6'h2e == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_46;
      end else if (6'h2d == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_45;
      end else if (6'h2c == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_44;
      end else if (6'h2b == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_43;
      end else if (6'h2a == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_42;
      end else if (6'h29 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_41;
      end else if (6'h28 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_40;
      end else if (6'h27 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_39;
      end else if (6'h26 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_38;
      end else if (6'h25 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_37;
      end else if (6'h24 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_36;
      end else if (6'h23 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_35;
      end else if (6'h22 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_34;
      end else if (6'h21 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_33;
      end else if (6'h20 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_32;
      end else if (6'h1f == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_31;
      end else if (6'h1e == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_30;
      end else if (6'h1d == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_29;
      end else if (6'h1c == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_28;
      end else if (6'h1b == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_27;
      end else if (6'h1a == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_26;
      end else if (6'h19 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_25;
      end else if (6'h18 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_24;
      end else if (6'h17 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_23;
      end else if (6'h16 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_22;
      end else if (6'h15 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_21;
      end else if (6'h14 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_20;
      end else if (6'h13 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_19;
      end else if (6'h12 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_18;
      end else if (6'h11 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_17;
      end else if (6'h10 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_16;
      end else if (6'hf == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_15;
      end else if (6'he == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_14;
      end else if (6'hd == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_13;
      end else if (6'hc == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_12;
      end else if (6'hb == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_11;
      end else if (6'ha == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_10;
      end else if (6'h9 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_9;
      end else if (6'h8 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_8;
      end else if (6'h7 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_7;
      end else if (6'h6 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_6;
      end else if (6'h5 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_5;
      end else if (6'h4 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_4;
      end else if (6'h3 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_3;
      end else if (6'h2 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_2;
      end else if (6'h1 == _T_969[5:0]) begin
        leftNeighb <= laggWindow_io_parallelOut_1;
      end else begin
        leftNeighb <= _GEN_655;
      end
    end else if (3'h7 == _T_972[2:0]) begin
      leftNeighb <= laggGuard_io_parallelOut_7;
    end else if (3'h6 == _T_972[2:0]) begin
      leftNeighb <= laggGuard_io_parallelOut_6;
    end else if (3'h5 == _T_972[2:0]) begin
      leftNeighb <= laggGuard_io_parallelOut_5;
    end else if (3'h4 == _T_972[2:0]) begin
      leftNeighb <= laggGuard_io_parallelOut_4;
    end else if (3'h3 == _T_972[2:0]) begin
      leftNeighb <= laggGuard_io_parallelOut_3;
    end else if (3'h2 == _T_972[2:0]) begin
      leftNeighb <= laggGuard_io_parallelOut_2;
    end else if (3'h1 == _T_972[2:0]) begin
      leftNeighb <= laggGuard_io_parallelOut_1;
    end else begin
      leftNeighb <= _GEN_719;
    end
    if (_T_967) begin
      rightNeighb <= leadWindow_io_parallelOut_0;
    end else begin
      rightNeighb <= leadGuard_io_parallelOut_0;
    end
    _T_985 <= initialInDone & _T_114;
    _T_986 <= io_out_ready;
    _T_993 <= initialInDone & _T_114;
    _T_994 <= io_out_ready;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3) begin
          $fwrite(32'h80000002,"Assertion failed: Number of window cells must be larger than number of sub cells\n    at CFARCoreWithASR.scala:20 assert(io.windowCells >= io.subCells.get, \"Number of window cells must be larger than number of sub cells\")\n"); // @[CFARCoreWithASR.scala 20:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3) begin
          $fatal; // @[CFARCoreWithASR.scala 20:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14) begin
          $fwrite(32'h80000002,"Assertion failed: FFT size must be larger than total number of shifting cells inside CFAR core\n    at CFARCoreWithASR.scala:38 assert(io.fftWin > 2.U * io.windowCells + 2.U * io.guardCells + 1.U, \"FFT size must be larger than total number of shifting cells inside CFAR core\")\n"); // @[CFARCoreWithASR.scala 38:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_14) begin
          $fatal; // @[CFARCoreWithASR.scala 38:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CFARCore(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input  [9:0]  io_fftWin,
  input  [15:0] io_thresholdScaler,
  input  [2:0]  io_divSum,
  input         io_peakGrouping,
  input  [1:0]  io_cfarMode,
  input  [6:0]  io_windowCells,
  input  [3:0]  io_guardCells,
  input  [6:0]  io_subCells,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_peak,
  output [15:0] io_out_bits_cut,
  output [15:0] io_out_bits_threshold,
  output        io_lastOut,
  output [8:0]  io_fftBin
);
  wire  cfarCore_clock; // @[CFARcore.scala 64:94]
  wire  cfarCore_reset; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_in_ready; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_in_valid; // @[CFARcore.scala 64:94]
  wire [15:0] cfarCore_io_in_bits; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_lastIn; // @[CFARcore.scala 64:94]
  wire [9:0] cfarCore_io_fftWin; // @[CFARcore.scala 64:94]
  wire [15:0] cfarCore_io_thresholdScaler; // @[CFARcore.scala 64:94]
  wire [2:0] cfarCore_io_divSum; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_peakGrouping; // @[CFARcore.scala 64:94]
  wire [1:0] cfarCore_io_cfarMode; // @[CFARcore.scala 64:94]
  wire [6:0] cfarCore_io_windowCells; // @[CFARcore.scala 64:94]
  wire [3:0] cfarCore_io_guardCells; // @[CFARcore.scala 64:94]
  wire [6:0] cfarCore_io_subCells; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_out_ready; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_out_valid; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_out_bits_peak; // @[CFARcore.scala 64:94]
  wire [15:0] cfarCore_io_out_bits_cut; // @[CFARcore.scala 64:94]
  wire [15:0] cfarCore_io_out_bits_threshold; // @[CFARcore.scala 64:94]
  wire  cfarCore_io_lastOut; // @[CFARcore.scala 64:94]
  wire [8:0] cfarCore_io_fftBin; // @[CFARcore.scala 64:94]
  CFARCoreWithASR cfarCore ( // @[CFARcore.scala 64:94]
    .clock(cfarCore_clock),
    .reset(cfarCore_reset),
    .io_in_ready(cfarCore_io_in_ready),
    .io_in_valid(cfarCore_io_in_valid),
    .io_in_bits(cfarCore_io_in_bits),
    .io_lastIn(cfarCore_io_lastIn),
    .io_fftWin(cfarCore_io_fftWin),
    .io_thresholdScaler(cfarCore_io_thresholdScaler),
    .io_divSum(cfarCore_io_divSum),
    .io_peakGrouping(cfarCore_io_peakGrouping),
    .io_cfarMode(cfarCore_io_cfarMode),
    .io_windowCells(cfarCore_io_windowCells),
    .io_guardCells(cfarCore_io_guardCells),
    .io_subCells(cfarCore_io_subCells),
    .io_out_ready(cfarCore_io_out_ready),
    .io_out_valid(cfarCore_io_out_valid),
    .io_out_bits_peak(cfarCore_io_out_bits_peak),
    .io_out_bits_cut(cfarCore_io_out_bits_cut),
    .io_out_bits_threshold(cfarCore_io_out_bits_threshold),
    .io_lastOut(cfarCore_io_lastOut),
    .io_fftBin(cfarCore_io_fftBin)
  );
  assign io_in_ready = cfarCore_io_in_ready; // @[CFARcore.scala 68:18]
  assign io_out_valid = cfarCore_io_out_valid; // @[CFARcore.scala 95:19]
  assign io_out_bits_peak = cfarCore_io_out_bits_peak; // @[CFARcore.scala 95:19]
  assign io_out_bits_cut = cfarCore_io_out_bits_cut; // @[CFARcore.scala 95:19]
  assign io_out_bits_threshold = cfarCore_io_out_bits_threshold; // @[CFARcore.scala 95:19]
  assign io_lastOut = cfarCore_io_lastOut; // @[CFARcore.scala 96:14]
  assign io_fftBin = cfarCore_io_fftBin; // @[CFARcore.scala 97:13]
  assign cfarCore_clock = clock;
  assign cfarCore_reset = reset;
  assign cfarCore_io_in_valid = io_in_valid; // @[CFARcore.scala 68:18]
  assign cfarCore_io_in_bits = io_in_bits; // @[CFARcore.scala 68:18]
  assign cfarCore_io_lastIn = io_lastIn; // @[CFARcore.scala 69:22]
  assign cfarCore_io_fftWin = io_fftWin; // @[CFARcore.scala 70:22]
  assign cfarCore_io_thresholdScaler = io_thresholdScaler; // @[CFARcore.scala 71:31]
  assign cfarCore_io_divSum = io_divSum; // @[CFARcore.scala 77:28]
  assign cfarCore_io_peakGrouping = io_peakGrouping; // @[CFARcore.scala 79:28]
  assign cfarCore_io_cfarMode = io_cfarMode; // @[CFARcore.scala 83:24]
  assign cfarCore_io_windowCells = io_windowCells; // @[CFARcore.scala 84:27]
  assign cfarCore_io_guardCells = io_guardCells; // @[CFARcore.scala 85:26]
  assign cfarCore_io_subCells = io_subCells; // @[CFARcore.scala 93:30]
  assign cfarCore_io_out_ready = io_out_ready; // @[CFARcore.scala 95:19]
endmodule
module AXI4CFARBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  input         auto_master_out_ready,
  output        auto_master_out_valid,
  output [47:0] auto_master_out_bits_data,
  output        auto_master_out_bits_last,
  output        auto_slave_in_ready,
  input         auto_slave_in_valid,
  input  [15:0] auto_slave_in_bits_data,
  input         auto_slave_in_bits_last
);
  wire  cfar_clock; // @[CFARDspBlock.scala 66:22]
  wire  cfar_reset; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_in_ready; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_in_valid; // @[CFARDspBlock.scala 66:22]
  wire [15:0] cfar_io_in_bits; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_lastIn; // @[CFARDspBlock.scala 66:22]
  wire [9:0] cfar_io_fftWin; // @[CFARDspBlock.scala 66:22]
  wire [15:0] cfar_io_thresholdScaler; // @[CFARDspBlock.scala 66:22]
  wire [2:0] cfar_io_divSum; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_peakGrouping; // @[CFARDspBlock.scala 66:22]
  wire [1:0] cfar_io_cfarMode; // @[CFARDspBlock.scala 66:22]
  wire [6:0] cfar_io_windowCells; // @[CFARDspBlock.scala 66:22]
  wire [3:0] cfar_io_guardCells; // @[CFARDspBlock.scala 66:22]
  wire [6:0] cfar_io_subCells; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_out_ready; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_out_valid; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_out_bits_peak; // @[CFARDspBlock.scala 66:22]
  wire [15:0] cfar_io_out_bits_cut; // @[CFARDspBlock.scala 66:22]
  wire [15:0] cfar_io_out_bits_threshold; // @[CFARDspBlock.scala 66:22]
  wire  cfar_io_lastOut; // @[CFARDspBlock.scala 66:22]
  wire [8:0] cfar_io_fftBin; // @[CFARDspBlock.scala 66:22]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [9:0] fftWin; // @[CFARDspBlock.scala 72:25]
  reg [31:0] _RAND_0;
  reg [15:0] thresholdScaler; // @[CFARDspBlock.scala 73:34]
  reg [31:0] _RAND_1;
  reg  peakGrouping; // @[CFARDspBlock.scala 74:31]
  reg [31:0] _RAND_2;
  reg [1:0] cfarMode; // @[CFARDspBlock.scala 75:27]
  reg [31:0] _RAND_3;
  reg [6:0] windowCells; // @[CFARDspBlock.scala 76:30]
  reg [31:0] _RAND_4;
  reg [3:0] guardCells; // @[CFARDspBlock.scala 77:29]
  reg [31:0] _RAND_5;
  reg [2:0] _T_6; // @[CFARDspBlock.scala 111:27]
  reg [31:0] _RAND_6;
  reg [6:0] subWindowSize; // @[CFARDspBlock.scala 118:34]
  reg [31:0] _RAND_7;
  wire [41:0] _T_11; // @[Cat.scala 29:58]
  wire  _T_13; // @[RegisterRouter.scala 40:39]
  wire  _T_14; // @[RegisterRouter.scala 40:26]
  wire  _T_15; // @[RegisterRouter.scala 42:29]
  wire  _T_58_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_22; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_312; // @[Cat.scala 29:58]
  wire [5:0] _T_62; // @[RegisterRouter.scala 59:16]
  wire  _T_74; // @[RegisterRouter.scala 59:16]
  wire  _T_16; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_25; // @[OneHot.scala 65:12]
  wire [1:0] _T_27; // @[Misc.scala 200:81]
  wire  _T_28; // @[Misc.scala 204:21]
  wire  _T_31; // @[Misc.scala 209:20]
  wire  _T_33; // @[Misc.scala 213:38]
  wire  _T_34; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 209:20]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 212:27]
  wire  _T_45; // @[Misc.scala 213:38]
  wire  _T_46; // @[Misc.scala 213:29]
  wire  _T_47; // @[Misc.scala 212:27]
  wire  _T_48; // @[Misc.scala 213:38]
  wire  _T_49; // @[Misc.scala 213:29]
  wire  _T_50; // @[Misc.scala 212:27]
  wire  _T_51; // @[Misc.scala 213:38]
  wire  _T_52; // @[Misc.scala 213:29]
  wire [3:0] _T_55; // @[Cat.scala 29:58]
  wire [3:0] _T_57; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_88; // @[Bitwise.scala 72:12]
  wire [7:0] _T_90; // @[Bitwise.scala 72:12]
  wire [7:0] _T_92; // @[Bitwise.scala 72:12]
  wire [7:0] _T_94; // @[Bitwise.scala 72:12]
  wire [31:0] _T_97; // @[Cat.scala 29:58]
  wire  _T_116; // @[RegisterRouter.scala 59:16]
  wire  _T_331; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_313; // @[OneHot.scala 58:35]
  wire  _T_378; // @[RegisterRouter.scala 59:16]
  wire  _T_380; // @[RegisterRouter.scala 59:16]
  wire  _T_381; // @[RegisterRouter.scala 59:16]
  wire  _T_123; // @[RegisterRouter.scala 59:16]
  wire  _T_139; // @[RegisterRouter.scala 59:16]
  wire  _T_405; // @[RegisterRouter.scala 59:16]
  wire  _T_406; // @[RegisterRouter.scala 59:16]
  wire  _T_146; // @[RegisterRouter.scala 59:16]
  wire  _T_162; // @[RegisterRouter.scala 59:16]
  wire  _T_385; // @[RegisterRouter.scala 59:16]
  wire  _T_386; // @[RegisterRouter.scala 59:16]
  wire  _T_169; // @[RegisterRouter.scala 59:16]
  wire  _T_185; // @[RegisterRouter.scala 59:16]
  wire  _T_410; // @[RegisterRouter.scala 59:16]
  wire  _T_411; // @[RegisterRouter.scala 59:16]
  wire  _T_192; // @[RegisterRouter.scala 59:16]
  wire  _T_390; // @[RegisterRouter.scala 59:16]
  wire  _T_391; // @[RegisterRouter.scala 59:16]
  wire  _T_215; // @[RegisterRouter.scala 59:16]
  wire  _T_231; // @[RegisterRouter.scala 59:16]
  wire  _T_415; // @[RegisterRouter.scala 59:16]
  wire  _T_416; // @[RegisterRouter.scala 59:16]
  wire  _T_238; // @[RegisterRouter.scala 59:16]
  wire  _T_254; // @[RegisterRouter.scala 59:16]
  wire  _T_395; // @[RegisterRouter.scala 59:16]
  wire  _T_396; // @[RegisterRouter.scala 59:16]
  wire  _T_261; // @[RegisterRouter.scala 59:16]
  wire  _T_400; // @[RegisterRouter.scala 59:16]
  wire  _T_401; // @[RegisterRouter.scala 59:16]
  wire  _T_284; // @[RegisterRouter.scala 59:16]
  wire  _GEN_41; // @[MuxLiteral.scala 48:10]
  wire  _GEN_42; // @[MuxLiteral.scala 48:10]
  wire  _GEN_43; // @[MuxLiteral.scala 48:10]
  wire  _GEN_44; // @[MuxLiteral.scala 48:10]
  wire  _GEN_45; // @[MuxLiteral.scala 48:10]
  wire  _GEN_46; // @[MuxLiteral.scala 48:10]
  wire  _GEN_47; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_523_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_49; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_523_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_50; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_523_3; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_51; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_523_4; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_52; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_523_5; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_53; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_523_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_54; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_523_7; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_55; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_525; // @[RegisterRouter.scala 59:16]
  wire  _T_526_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_526_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_529; // @[RegisterRouter.scala 65:29]
  CFARCore cfar ( // @[CFARDspBlock.scala 66:22]
    .clock(cfar_clock),
    .reset(cfar_reset),
    .io_in_ready(cfar_io_in_ready),
    .io_in_valid(cfar_io_in_valid),
    .io_in_bits(cfar_io_in_bits),
    .io_lastIn(cfar_io_lastIn),
    .io_fftWin(cfar_io_fftWin),
    .io_thresholdScaler(cfar_io_thresholdScaler),
    .io_divSum(cfar_io_divSum),
    .io_peakGrouping(cfar_io_peakGrouping),
    .io_cfarMode(cfar_io_cfarMode),
    .io_windowCells(cfar_io_windowCells),
    .io_guardCells(cfar_io_guardCells),
    .io_subCells(cfar_io_subCells),
    .io_out_ready(cfar_io_out_ready),
    .io_out_valid(cfar_io_out_valid),
    .io_out_bits_peak(cfar_io_out_bits_peak),
    .io_out_bits_cut(cfar_io_out_bits_cut),
    .io_out_bits_threshold(cfar_io_out_bits_threshold),
    .io_lastOut(cfar_io_lastOut),
    .io_fftBin(cfar_io_fftBin)
  );
  Queue_1 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_11 = {cfar_io_out_bits_threshold,cfar_io_out_bits_cut,cfar_io_fftBin,cfar_io_out_bits_peak}; // @[Cat.scala 29:58]
  assign _T_13 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_14 = auto_mem_in_ar_valid | _T_13; // @[RegisterRouter.scala 40:26]
  assign _T_15 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_58_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_22 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_312 = {_T_22[4],_T_22[3],_T_22[2]}; // @[Cat.scala 29:58]
  assign _T_62 = _T_22[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  assign _T_74 = _T_62 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_16 = _T_58_ready & _T_15; // @[RegisterRouter.scala 42:26]
  assign _T_25 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_27 = _T_25 | 2'h1; // @[Misc.scala 200:81]
  assign _T_28 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_31 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_33 = _T_27[1] & _T_31; // @[Misc.scala 213:38]
  assign _T_34 = _T_28 | _T_33; // @[Misc.scala 213:29]
  assign _T_36 = _T_27[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_37 = _T_28 | _T_36; // @[Misc.scala 213:29]
  assign _T_40 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_41 = _T_31 & _T_40; // @[Misc.scala 212:27]
  assign _T_42 = _T_27[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_34 | _T_42; // @[Misc.scala 213:29]
  assign _T_44 = _T_31 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_45 = _T_27[0] & _T_44; // @[Misc.scala 213:38]
  assign _T_46 = _T_34 | _T_45; // @[Misc.scala 213:29]
  assign _T_47 = auto_mem_in_ar_bits_addr[1] & _T_40; // @[Misc.scala 212:27]
  assign _T_48 = _T_27[0] & _T_47; // @[Misc.scala 213:38]
  assign _T_49 = _T_37 | _T_48; // @[Misc.scala 213:29]
  assign _T_50 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_51 = _T_27[0] & _T_50; // @[Misc.scala 213:38]
  assign _T_52 = _T_37 | _T_51; // @[Misc.scala 213:29]
  assign _T_55 = {_T_52,_T_49,_T_46,_T_43}; // @[Cat.scala 29:58]
  assign _T_57 = auto_mem_in_ar_valid ? _T_55 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_88 = _T_57[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_90 = _T_57[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_92 = _T_57[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_94 = _T_57[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_97 = {_T_94,_T_92,_T_90,_T_88}; // @[Cat.scala 29:58]
  assign _T_116 = _T_97[9:0] == 10'h3ff; // @[RegisterRouter.scala 59:16]
  assign _T_331 = _T_14 & _T_58_ready; // @[RegisterRouter.scala 59:16]
  assign _T_313 = 8'h1 << _T_312; // @[OneHot.scala 58:35]
  assign _T_378 = _T_331 & _T_15; // @[RegisterRouter.scala 59:16]
  assign _T_380 = _T_378 & _T_313[0]; // @[RegisterRouter.scala 59:16]
  assign _T_381 = _T_380 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_123 = _T_381 & _T_116; // @[RegisterRouter.scala 59:16]
  assign _T_139 = _T_97[3:0] == 4'hf; // @[RegisterRouter.scala 59:16]
  assign _T_405 = _T_378 & _T_313[5]; // @[RegisterRouter.scala 59:16]
  assign _T_406 = _T_405 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_146 = _T_406 & _T_139; // @[RegisterRouter.scala 59:16]
  assign _T_162 = _T_97[15:0] == 16'hffff; // @[RegisterRouter.scala 59:16]
  assign _T_385 = _T_378 & _T_313[1]; // @[RegisterRouter.scala 59:16]
  assign _T_386 = _T_385 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_169 = _T_386 & _T_162; // @[RegisterRouter.scala 59:16]
  assign _T_185 = _T_97[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_410 = _T_378 & _T_313[6]; // @[RegisterRouter.scala 59:16]
  assign _T_411 = _T_410 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_192 = _T_411 & _T_185; // @[RegisterRouter.scala 59:16]
  assign _T_390 = _T_378 & _T_313[2]; // @[RegisterRouter.scala 59:16]
  assign _T_391 = _T_390 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_215 = _T_391 & _T_97[0]; // @[RegisterRouter.scala 59:16]
  assign _T_231 = _T_97[6:0] == 7'h7f; // @[RegisterRouter.scala 59:16]
  assign _T_415 = _T_378 & _T_313[7]; // @[RegisterRouter.scala 59:16]
  assign _T_416 = _T_415 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_238 = _T_416 & _T_231; // @[RegisterRouter.scala 59:16]
  assign _T_254 = _T_97[1:0] == 2'h3; // @[RegisterRouter.scala 59:16]
  assign _T_395 = _T_378 & _T_313[3]; // @[RegisterRouter.scala 59:16]
  assign _T_396 = _T_395 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_261 = _T_396 & _T_254; // @[RegisterRouter.scala 59:16]
  assign _T_400 = _T_378 & _T_313[4]; // @[RegisterRouter.scala 59:16]
  assign _T_401 = _T_400 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_284 = _T_401 & _T_231; // @[RegisterRouter.scala 59:16]
  assign _GEN_41 = 3'h1 == _T_312 ? _T_74 : _T_74; // @[MuxLiteral.scala 48:10]
  assign _GEN_42 = 3'h2 == _T_312 ? _T_74 : _GEN_41; // @[MuxLiteral.scala 48:10]
  assign _GEN_43 = 3'h3 == _T_312 ? _T_74 : _GEN_42; // @[MuxLiteral.scala 48:10]
  assign _GEN_44 = 3'h4 == _T_312 ? _T_74 : _GEN_43; // @[MuxLiteral.scala 48:10]
  assign _GEN_45 = 3'h5 == _T_312 ? _T_74 : _GEN_44; // @[MuxLiteral.scala 48:10]
  assign _GEN_46 = 3'h6 == _T_312 ? _T_74 : _GEN_45; // @[MuxLiteral.scala 48:10]
  assign _GEN_47 = 3'h7 == _T_312 ? _T_74 : _GEN_46; // @[MuxLiteral.scala 48:10]
  assign _T_523_0 = {{6'd0}, fftWin}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_49 = 3'h1 == _T_312 ? thresholdScaler : _T_523_0; // @[MuxLiteral.scala 48:10]
  assign _T_523_2 = {{15'd0}, peakGrouping}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_50 = 3'h2 == _T_312 ? _T_523_2 : _GEN_49; // @[MuxLiteral.scala 48:10]
  assign _T_523_3 = {{14'd0}, cfarMode}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_51 = 3'h3 == _T_312 ? _T_523_3 : _GEN_50; // @[MuxLiteral.scala 48:10]
  assign _T_523_4 = {{9'd0}, windowCells}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_52 = 3'h4 == _T_312 ? _T_523_4 : _GEN_51; // @[MuxLiteral.scala 48:10]
  assign _T_523_5 = {{12'd0}, guardCells}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_53 = 3'h5 == _T_312 ? _T_523_5 : _GEN_52; // @[MuxLiteral.scala 48:10]
  assign _T_523_6 = {{13'd0}, _T_6}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_54 = 3'h6 == _T_312 ? _T_523_6 : _GEN_53; // @[MuxLiteral.scala 48:10]
  assign _T_523_7 = {{9'd0}, subWindowSize}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_55 = 3'h7 == _T_312 ? _T_523_7 : _GEN_54; // @[MuxLiteral.scala 48:10]
  assign _T_525 = _GEN_47 ? _GEN_55 : 16'h0; // @[RegisterRouter.scala 59:16]
  assign _T_526_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_526_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_529 = ~_T_526_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_16 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_16 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_526_valid & _T_529; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_526_valid & _T_526_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_master_out_valid = cfar_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_data = {{6'd0}, _T_11}; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_last = cfar_io_lastOut; // @[LazyModule.scala 173:49]
  assign auto_slave_in_ready = cfar_io_in_ready; // @[LazyModule.scala 173:31]
  assign cfar_clock = clock;
  assign cfar_reset = reset;
  assign cfar_io_in_valid = auto_slave_in_valid; // @[CFARDspBlock.scala 97:22]
  assign cfar_io_in_bits = auto_slave_in_bits_data; // @[CFARDspBlock.scala 98:21]
  assign cfar_io_lastIn = auto_slave_in_bits_last; // @[CFARDspBlock.scala 135:25]
  assign cfar_io_fftWin = fftWin; // @[CFARDspBlock.scala 100:20]
  assign cfar_io_thresholdScaler = thresholdScaler; // @[CFARDspBlock.scala 101:29]
  assign cfar_io_divSum = _T_6; // @[CFARDspBlock.scala 112:26]
  assign cfar_io_peakGrouping = peakGrouping; // @[CFARDspBlock.scala 124:26]
  assign cfar_io_cfarMode = cfarMode; // @[CFARDspBlock.scala 132:25]
  assign cfar_io_windowCells = windowCells; // @[CFARDspBlock.scala 133:25]
  assign cfar_io_guardCells = guardCells; // @[CFARDspBlock.scala 134:25]
  assign cfar_io_subCells = subWindowSize; // @[CFARDspBlock.scala 122:28]
  assign cfar_io_out_ready = auto_master_out_ready; // @[CFARDspBlock.scala 162:24]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_13; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{16'd0}, _T_525}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_526_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fftWin = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  thresholdScaler = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  peakGrouping = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cfarMode = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  windowCells = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  guardCells = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  subWindowSize = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fftWin <= 10'h200;
    end else if (_T_123) begin
      fftWin <= auto_mem_in_w_bits_data[9:0];
    end
    if (reset) begin
      thresholdScaler <= 16'h0;
    end else if (_T_169) begin
      thresholdScaler <= auto_mem_in_w_bits_data[15:0];
    end
    if (reset) begin
      peakGrouping <= 1'h0;
    end else if (_T_215) begin
      peakGrouping <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      cfarMode <= 2'h0;
    end else if (_T_261) begin
      cfarMode <= auto_mem_in_w_bits_data[1:0];
    end
    if (reset) begin
      windowCells <= 7'h40;
    end else if (_T_284) begin
      windowCells <= auto_mem_in_w_bits_data[6:0];
    end
    if (reset) begin
      guardCells <= 4'h8;
    end else if (_T_146) begin
      guardCells <= auto_mem_in_w_bits_data[3:0];
    end
    if (reset) begin
      _T_6 <= 3'h0;
    end else if (_T_192) begin
      _T_6 <= auto_mem_in_w_bits_data[2:0];
    end
    if (reset) begin
      subWindowSize <= 7'h0;
    end else if (_T_238) begin
      subWindowSize <= auto_mem_in_w_bits_data[6:0];
    end
  end
endmodule
module AXI4StreamWidthAdapater_1_to_3(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [47:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [15:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [1:0] _T_4; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_0;
  wire  _T_5; // @[AXI4StreamWidthAdapter.scala 159:14]
  wire  _T_6; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_7; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_8; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir0; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_10; // @[AXI4StreamWidthAdapter.scala 167:22]
  reg [31:0] _RAND_1;
  wire  _T_12; // @[AXI4StreamWidthAdapter.scala 168:38]
  wire [2:0] _T_13; // @[AXI4StreamWidthAdapter.scala 168:60]
  wire [2:0] _T_14; // @[AXI4StreamWidthAdapter.scala 168:33]
  wire [2:0] _GEN_1; // @[AXI4StreamWidthAdapter.scala 168:21]
  wire  ir1; // @[AXI4StreamWidthAdapter.scala 170:60]
  reg [1:0] _T_19; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_2;
  wire  _T_21; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_22; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_23; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_2; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir2; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_26; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_3;
  wire  _T_28; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_29; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_30; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_3; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir3; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_33; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_4;
  wire  _T_35; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_36; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_37; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir4; // @[AXI4StreamWidthAdapter.scala 163:34]
  wire  _T_55; // @[AXI4StreamWidthAdapter.scala 46:16]
  wire  _T_57; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_58; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_59; // @[AXI4StreamWidthAdapter.scala 47:16]
  wire  _T_61; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_62; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_63; // @[AXI4StreamWidthAdapter.scala 48:16]
  wire  _T_65; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_67; // @[AXI4StreamWidthAdapter.scala 49:16]
  wire  _T_69; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire  _T_70; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire [15:0] _GEN_6; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign _T_5 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 159:14]
  assign _T_6 = _T_4 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_7 = _T_4 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_8 = _T_6 ? 3'h0 : _T_7; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_0 = _T_5 ? _T_8 : {{1'd0}, _T_4}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir0 = _T_6 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_12 = _T_10 == 2'h2; // @[AXI4StreamWidthAdapter.scala 168:38]
  assign _T_13 = _T_10 + 2'h1; // @[AXI4StreamWidthAdapter.scala 168:60]
  assign _T_14 = _T_12 ? 3'h0 : _T_13; // @[AXI4StreamWidthAdapter.scala 168:33]
  assign _GEN_1 = _T_5 ? _T_14 : {{1'd0}, _T_10}; // @[AXI4StreamWidthAdapter.scala 168:21]
  assign ir1 = _T_12 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 170:60]
  assign _T_21 = _T_19 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_22 = _T_19 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_23 = _T_21 ? 3'h0 : _T_22; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_2 = _T_5 ? _T_23 : {{1'd0}, _T_19}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir2 = _T_21 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_28 = _T_26 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_29 = _T_26 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_30 = _T_28 ? 3'h0 : _T_29; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_3 = _T_5 ? _T_30 : {{1'd0}, _T_26}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir3 = _T_28 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_35 = _T_33 == 2'h2; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_36 = _T_33 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_37 = _T_35 ? 3'h0 : _T_36; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_4 = _T_5 ? _T_37 : {{1'd0}, _T_33}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir4 = _T_35 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_55 = ir0 == ir1; // @[AXI4StreamWidthAdapter.scala 46:16]
  assign _T_57 = _T_55 | reset; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign _T_58 = ~_T_57; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign _T_59 = ir0 == ir2; // @[AXI4StreamWidthAdapter.scala 47:16]
  assign _T_61 = _T_59 | reset; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign _T_62 = ~_T_61; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign _T_63 = ir0 == ir3; // @[AXI4StreamWidthAdapter.scala 48:16]
  assign _T_65 = _T_63 | reset; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign _T_66 = ~_T_65; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign _T_67 = ir0 == ir4; // @[AXI4StreamWidthAdapter.scala 49:16]
  assign _T_69 = _T_67 | reset; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign _T_70 = ~_T_69; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign _GEN_6 = 2'h1 == _T_4 ? auto_in_bits_data[31:16] : auto_in_bits_data[15:0]; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign auto_in_ready = _T_6 & auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = 2'h2 == _T_4 ? auto_in_bits_data[47:32] : _GEN_6; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last & _T_12; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_19 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_33 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_4 <= 2'h0;
    end else begin
      _T_4 <= _GEN_0[1:0];
    end
    if (reset) begin
      _T_10 <= 2'h0;
    end else begin
      _T_10 <= _GEN_1[1:0];
    end
    if (reset) begin
      _T_19 <= 2'h0;
    end else begin
      _T_19 <= _GEN_2[1:0];
    end
    if (reset) begin
      _T_26 <= 2'h0;
    end else begin
      _T_26 <= _GEN_3[1:0];
    end
    if (reset) begin
      _T_33 <= 2'h0;
    end else begin
      _T_33 <= _GEN_4[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_58) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:46 assert(ir0 === ir1)\n"); // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_58) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_62) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:47 assert(ir0 === ir2)\n"); // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_62) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_66) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:48 assert(ir0 === ir3)\n"); // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_66) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_70) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:49 assert(ir0 === ir4)\n"); // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_70) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_8 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_9(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [15:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [15:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [15:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [15:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [15:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_9 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_11(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [47:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [47:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [47:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [63:0] _RAND_0;
  wire [47:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [47:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[47:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_3(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [47:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [47:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [47:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [47:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_11 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module QueueCompatibility(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits
);
  reg [2:0] _T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [2:0] _T__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [2:0] _T__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _GEN_9; // @[Decoupled.scala 240:27]
  wire  _GEN_12; // @[Decoupled.scala 237:18]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _GEN_11; // @[Decoupled.scala 237:18]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire  _T_16; // @[Decoupled.scala 231:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = _T_4 ? _GEN_9 : _T_6;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_12 = _T_4 ? _GEN_9 : _T_6; // @[Decoupled.scala 237:18]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_11 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_15 = _GEN_12 != _GEN_11; // @[Decoupled.scala 227:16]
  assign _T_16 = ~_T_4; // @[Decoupled.scala 231:19]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = _T_4 ? io_enq_bits : _T__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_12) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_11) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module AXI4Xbar(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_2_aw_ready,
  output        auto_out_2_aw_valid,
  output        auto_out_2_aw_bits_id,
  output [29:0] auto_out_2_aw_bits_addr,
  input         auto_out_2_w_ready,
  output        auto_out_2_w_valid,
  output [31:0] auto_out_2_w_bits_data,
  output [3:0]  auto_out_2_w_bits_strb,
  output        auto_out_2_b_ready,
  input         auto_out_2_b_valid,
  input         auto_out_2_b_bits_id,
  input         auto_out_2_ar_ready,
  output        auto_out_2_ar_valid,
  output        auto_out_2_ar_bits_id,
  output [29:0] auto_out_2_ar_bits_addr,
  output [2:0]  auto_out_2_ar_bits_size,
  output        auto_out_2_r_ready,
  input         auto_out_2_r_valid,
  input         auto_out_2_r_bits_id,
  input  [31:0] auto_out_2_r_bits_data,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output        auto_out_0_aw_bits_id,
  output [29:0] auto_out_0_aw_bits_addr,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid,
  input         auto_out_0_b_bits_id,
  input         auto_out_0_ar_ready,
  output        auto_out_0_ar_valid,
  output        auto_out_0_ar_bits_id,
  output [29:0] auto_out_0_ar_bits_addr,
  output        auto_out_0_r_ready,
  input         auto_out_0_r_valid,
  input         auto_out_0_r_bits_id,
  input  [31:0] auto_out_0_r_bits_data
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [2:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [2:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1; // @[Parameters.scala 137:49]
  wire [30:0] _T_3; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5; // @[Parameters.scala 137:31]
  wire [30:0] _T_6; // @[Parameters.scala 137:49]
  wire [30:0] _T_8; // @[Parameters.scala 137:52]
  wire  requestARIO_0_1; // @[Parameters.scala 137:67]
  wire [29:0] _T_10; // @[Parameters.scala 137:31]
  wire [30:0] _T_11; // @[Parameters.scala 137:49]
  wire [30:0] _T_13; // @[Parameters.scala 137:52]
  wire  requestARIO_0_2; // @[Parameters.scala 137:67]
  wire [30:0] _T_16; // @[Parameters.scala 137:49]
  wire [30:0] _T_18; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_20; // @[Parameters.scala 137:31]
  wire [30:0] _T_21; // @[Parameters.scala 137:49]
  wire [30:0] _T_23; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_1; // @[Parameters.scala 137:67]
  wire [29:0] _T_25; // @[Parameters.scala 137:31]
  wire [30:0] _T_26; // @[Parameters.scala 137:49]
  wire [30:0] _T_28; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_2; // @[Parameters.scala 137:67]
  wire  requestROI_0_0; // @[Parameters.scala 47:9]
  wire  requestROI_1_0; // @[Parameters.scala 47:9]
  wire  requestROI_2_0; // @[Parameters.scala 47:9]
  wire  requestBOI_0_0; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0; // @[Parameters.scala 47:9]
  wire  requestBOI_2_0; // @[Parameters.scala 47:9]
  wire [1:0] _T_30; // @[Xbar.scala 64:75]
  wire [2:0] _T_31; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1; // @[Xbar.scala 65:73]
  wire  requestWIO_0_2; // @[Xbar.scala 65:73]
  wire [2:0] _T_39; // @[Xbar.scala 93:45]
  wire [1:0] _GEN_22; // @[OneHot.scala 32:28]
  wire [1:0] _T_43; // @[OneHot.scala 32:28]
  wire [1:0] _T_45; // @[Cat.scala 29:58]
  wire [1:0] _GEN_23; // @[OneHot.scala 32:28]
  wire [1:0] _T_51; // @[OneHot.scala 32:28]
  wire [1:0] _T_53; // @[Cat.scala 29:58]
  wire  _T_132; // @[Mux.scala 27:72]
  wire  _T_133; // @[Mux.scala 27:72]
  wire  _T_135; // @[Mux.scala 27:72]
  wire  _T_134; // @[Mux.scala 27:72]
  wire  in_0_ar_ready; // @[Mux.scala 27:72]
  reg [2:0] _T_59; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_78; // @[Xbar.scala 112:22]
  reg [1:0] _T_60; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_77; // @[Xbar.scala 111:75]
  wire  _T_79; // @[Xbar.scala 112:34]
  wire  _T_80; // @[Xbar.scala 112:80]
  wire  _T_82; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready; // @[Xbar.scala 130:45]
  wire  _T_54; // @[Decoupled.scala 40:37]
  reg  _T_302; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_159; // @[Xbar.scala 222:40]
  wire  _T_161; // @[Xbar.scala 222:40]
  wire  _T_303; // @[Xbar.scala 246:36]
  wire  _T_163; // @[Xbar.scala 222:40]
  wire  _T_304; // @[Xbar.scala 246:36]
  reg  _T_373_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_380; // @[Mux.scala 27:72]
  reg  _T_373_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_4;
  wire  _T_381; // @[Mux.scala 27:72]
  wire  _T_383; // @[Mux.scala 27:72]
  reg  _T_373_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_5;
  wire  _T_382; // @[Mux.scala 27:72]
  wire  _T_384; // @[Mux.scala 27:72]
  wire  in_0_r_valid; // @[Xbar.scala 278:22]
  wire  _T_56; // @[Decoupled.scala 40:37]
  wire [2:0] _T_306; // @[Cat.scala 29:58]
  reg [2:0] _T_313; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_6;
  wire [2:0] _T_314; // @[Arbiter.scala 21:30]
  wire [2:0] _T_315; // @[Arbiter.scala 21:28]
  wire [5:0] _T_316; // @[Cat.scala 29:58]
  wire [5:0] _GEN_24; // @[package.scala 208:43]
  wire [5:0] _T_318; // @[package.scala 208:43]
  wire [5:0] _GEN_25; // @[package.scala 208:43]
  wire [5:0] _T_320; // @[package.scala 208:43]
  wire [5:0] _T_323; // @[Arbiter.scala 22:66]
  wire [5:0] _GEN_26; // @[Arbiter.scala 22:58]
  wire [5:0] _T_324; // @[Arbiter.scala 22:58]
  wire [2:0] _T_327; // @[Arbiter.scala 23:39]
  wire [2:0] _T_328; // @[Arbiter.scala 23:18]
  wire  _T_344; // @[Xbar.scala 250:63]
  wire  _T_374_0; // @[Xbar.scala 262:23]
  wire [35:0] _T_389; // @[Mux.scala 27:72]
  wire [35:0] _T_390; // @[Mux.scala 27:72]
  wire  _T_345; // @[Xbar.scala 250:63]
  wire  _T_374_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_393; // @[Mux.scala 27:72]
  wire [35:0] _T_394; // @[Mux.scala 27:72]
  wire [35:0] _T_399; // @[Mux.scala 27:72]
  wire  _T_346; // @[Xbar.scala 250:63]
  wire  _T_374_2; // @[Xbar.scala 262:23]
  wire [35:0] _T_397; // @[Mux.scala 27:72]
  wire [35:0] _T_398; // @[Mux.scala 27:72]
  wire [35:0] _T_400; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last; // @[Mux.scala 27:72]
  wire  _T_58; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_27; // @[Xbar.scala 106:30]
  wire [2:0] _T_62; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_28; // @[Xbar.scala 106:48]
  wire [2:0] _T_64; // @[Xbar.scala 106:48]
  wire  _T_65; // @[Xbar.scala 107:23]
  wire  _T_66; // @[Xbar.scala 107:43]
  wire  _T_67; // @[Xbar.scala 107:34]
  wire  _T_69; // @[Xbar.scala 107:22]
  wire  _T_70; // @[Xbar.scala 107:22]
  wire  _T_71; // @[Xbar.scala 108:23]
  wire  _T_73; // @[Xbar.scala 108:34]
  wire  _T_75; // @[Xbar.scala 108:22]
  wire  _T_76; // @[Xbar.scala 108:22]
  wire  _T_142; // @[Mux.scala 27:72]
  wire  _T_143; // @[Mux.scala 27:72]
  wire  _T_145; // @[Mux.scala 27:72]
  wire  _T_144; // @[Mux.scala 27:72]
  wire  in_0_aw_ready; // @[Mux.scala 27:72]
  reg  _T_113; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_7;
  wire  _T_117; // @[Xbar.scala 139:57]
  wire  _T_118; // @[Xbar.scala 139:45]
  reg [2:0] _T_87; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_8;
  wire  _T_106; // @[Xbar.scala 112:22]
  reg [1:0] _T_88; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_9;
  wire  _T_105; // @[Xbar.scala 111:75]
  wire  _T_107; // @[Xbar.scala 112:34]
  wire  _T_108; // @[Xbar.scala 112:80]
  wire  _T_110; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready; // @[Xbar.scala 139:82]
  wire  _T_83; // @[Decoupled.scala 40:37]
  reg  _T_407; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_10;
  wire  _T_165; // @[Xbar.scala 222:40]
  wire  _T_167; // @[Xbar.scala 222:40]
  wire  _T_408; // @[Xbar.scala 246:36]
  wire  _T_169; // @[Xbar.scala 222:40]
  wire  _T_409; // @[Xbar.scala 246:36]
  reg  _T_478_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_11;
  wire  _T_485; // @[Mux.scala 27:72]
  reg  _T_478_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_12;
  wire  _T_486; // @[Mux.scala 27:72]
  wire  _T_488; // @[Mux.scala 27:72]
  reg  _T_478_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_13;
  wire  _T_487; // @[Mux.scala 27:72]
  wire  _T_489; // @[Mux.scala 27:72]
  wire  in_0_b_valid; // @[Xbar.scala 278:22]
  wire  _T_85; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_29; // @[Xbar.scala 106:30]
  wire [2:0] _T_90; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_30; // @[Xbar.scala 106:48]
  wire [2:0] _T_92; // @[Xbar.scala 106:48]
  wire  _T_93; // @[Xbar.scala 107:23]
  wire  _T_94; // @[Xbar.scala 107:43]
  wire  _T_95; // @[Xbar.scala 107:34]
  wire  _T_97; // @[Xbar.scala 107:22]
  wire  _T_98; // @[Xbar.scala 107:22]
  wire  _T_99; // @[Xbar.scala 108:23]
  wire  _T_101; // @[Xbar.scala 108:34]
  wire  _T_103; // @[Xbar.scala 108:22]
  wire  _T_104; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid; // @[Xbar.scala 129:45]
  wire  _T_115; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid; // @[Xbar.scala 138:82]
  wire  _T_120; // @[Xbar.scala 140:54]
  wire  _T_122; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[Xbar.scala 141:38]
  wire  _T_123; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid; // @[Xbar.scala 145:43]
  wire  _T_152; // @[Mux.scala 27:72]
  wire  _T_153; // @[Mux.scala 27:72]
  wire  _T_155; // @[Mux.scala 27:72]
  wire  _T_154; // @[Mux.scala 27:72]
  wire  in_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_126; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid; // @[Xbar.scala 222:40]
  wire  out_2_ar_valid; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid; // @[Xbar.scala 222:40]
  wire  out_2_aw_valid; // @[Xbar.scala 222:40]
  wire  _T_176; // @[Xbar.scala 256:60]
  wire  _T_182; // @[Xbar.scala 258:23]
  wire  _T_184; // @[Xbar.scala 258:12]
  wire  _T_185; // @[Xbar.scala 258:12]
  wire  _T_197; // @[Xbar.scala 256:60]
  wire  _T_203; // @[Xbar.scala 258:23]
  wire  _T_205; // @[Xbar.scala 258:12]
  wire  _T_206; // @[Xbar.scala 258:12]
  wire  _T_220; // @[Xbar.scala 256:60]
  wire  _T_226; // @[Xbar.scala 258:23]
  wire  _T_228; // @[Xbar.scala 258:12]
  wire  _T_229; // @[Xbar.scala 258:12]
  wire  _T_241; // @[Xbar.scala 256:60]
  wire  _T_247; // @[Xbar.scala 258:23]
  wire  _T_249; // @[Xbar.scala 258:12]
  wire  _T_250; // @[Xbar.scala 258:12]
  wire  _T_264; // @[Xbar.scala 256:60]
  wire  _T_270; // @[Xbar.scala 258:23]
  wire  _T_272; // @[Xbar.scala 258:12]
  wire  _T_273; // @[Xbar.scala 258:12]
  wire  _T_285; // @[Xbar.scala 256:60]
  wire  _T_291; // @[Xbar.scala 258:23]
  wire  _T_293; // @[Xbar.scala 258:12]
  wire  _T_294; // @[Xbar.scala 258:12]
  wire  _T_329; // @[Arbiter.scala 24:27]
  wire  _T_330; // @[Arbiter.scala 24:18]
  wire [2:0] _T_331; // @[Arbiter.scala 25:29]
  wire [3:0] _T_332; // @[package.scala 199:48]
  wire [2:0] _T_334; // @[package.scala 199:43]
  wire [4:0] _T_335; // @[package.scala 199:48]
  wire [2:0] _T_337; // @[package.scala 199:43]
  wire  _T_349; // @[Xbar.scala 255:50]
  wire  _T_350; // @[Xbar.scala 255:50]
  wire  _T_352; // @[Xbar.scala 256:60]
  wire  _T_355; // @[Xbar.scala 256:60]
  wire  _T_356; // @[Xbar.scala 256:57]
  wire  _T_357; // @[Xbar.scala 256:54]
  wire  _T_358; // @[Xbar.scala 256:60]
  wire  _T_359; // @[Xbar.scala 256:57]
  wire  _T_361; // @[Xbar.scala 256:75]
  wire  _T_363; // @[Xbar.scala 256:11]
  wire  _T_364; // @[Xbar.scala 256:11]
  wire  _T_365; // @[Xbar.scala 258:13]
  wire  _T_368; // @[Xbar.scala 258:23]
  wire  _T_370; // @[Xbar.scala 258:12]
  wire  _T_371; // @[Xbar.scala 258:12]
  wire  _GEN_17; // @[Xbar.scala 266:21]
  wire  _GEN_18; // @[Xbar.scala 267:24]
  wire  _T_376_0; // @[Xbar.scala 270:24]
  wire  _T_376_1; // @[Xbar.scala 270:24]
  wire  _T_376_2; // @[Xbar.scala 270:24]
  wire [2:0] _T_411; // @[Cat.scala 29:58]
  reg [2:0] _T_418; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_14;
  wire [2:0] _T_419; // @[Arbiter.scala 21:30]
  wire [2:0] _T_420; // @[Arbiter.scala 21:28]
  wire [5:0] _T_421; // @[Cat.scala 29:58]
  wire [5:0] _GEN_31; // @[package.scala 208:43]
  wire [5:0] _T_423; // @[package.scala 208:43]
  wire [5:0] _GEN_32; // @[package.scala 208:43]
  wire [5:0] _T_425; // @[package.scala 208:43]
  wire [5:0] _T_428; // @[Arbiter.scala 22:66]
  wire [5:0] _GEN_33; // @[Arbiter.scala 22:58]
  wire [5:0] _T_429; // @[Arbiter.scala 22:58]
  wire [2:0] _T_432; // @[Arbiter.scala 23:39]
  wire [2:0] _T_433; // @[Arbiter.scala 23:18]
  wire  _T_434; // @[Arbiter.scala 24:27]
  wire  _T_435; // @[Arbiter.scala 24:18]
  wire [2:0] _T_436; // @[Arbiter.scala 25:29]
  wire [3:0] _T_437; // @[package.scala 199:48]
  wire [2:0] _T_439; // @[package.scala 199:43]
  wire [4:0] _T_440; // @[package.scala 199:48]
  wire [2:0] _T_442; // @[package.scala 199:43]
  wire  _T_449; // @[Xbar.scala 250:63]
  wire  _T_450; // @[Xbar.scala 250:63]
  wire  _T_451; // @[Xbar.scala 250:63]
  wire  _T_454; // @[Xbar.scala 255:50]
  wire  _T_455; // @[Xbar.scala 255:50]
  wire  _T_457; // @[Xbar.scala 256:60]
  wire  _T_460; // @[Xbar.scala 256:60]
  wire  _T_461; // @[Xbar.scala 256:57]
  wire  _T_462; // @[Xbar.scala 256:54]
  wire  _T_463; // @[Xbar.scala 256:60]
  wire  _T_464; // @[Xbar.scala 256:57]
  wire  _T_466; // @[Xbar.scala 256:75]
  wire  _T_468; // @[Xbar.scala 256:11]
  wire  _T_469; // @[Xbar.scala 256:11]
  wire  _T_470; // @[Xbar.scala 258:13]
  wire  _T_473; // @[Xbar.scala 258:23]
  wire  _T_475; // @[Xbar.scala 258:12]
  wire  _T_476; // @[Xbar.scala 258:12]
  wire  _T_479_0; // @[Xbar.scala 262:23]
  wire  _T_479_1; // @[Xbar.scala 262:23]
  wire  _T_479_2; // @[Xbar.scala 262:23]
  wire  _GEN_20; // @[Xbar.scala 266:21]
  wire  _GEN_21; // @[Xbar.scala 267:24]
  wire  _T_481_0; // @[Xbar.scala 270:24]
  wire  _T_481_1; // @[Xbar.scala 270:24]
  wire  _T_481_2; // @[Xbar.scala 270:24]
  wire [2:0] _T_492; // @[Mux.scala 27:72]
  wire [2:0] _T_493; // @[Mux.scala 27:72]
  wire [2:0] _T_494; // @[Mux.scala 27:72]
  wire [2:0] _T_495; // @[Mux.scala 27:72]
  wire [2:0] _T_496; // @[Mux.scala 27:72]
  wire [2:0] _T_497; // @[Mux.scala 27:72]
  wire [2:0] _T_498; // @[Mux.scala 27:72]
  wire [2:0] _T_499; // @[Mux.scala 27:72]
  QueueCompatibility awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_3 = $signed(_T_1) & 31'sh300; // @[Parameters.scala 137:52]
  assign requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_5 = auto_in_ar_bits_addr ^ 30'h100; // @[Parameters.scala 137:31]
  assign _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  assign _T_8 = $signed(_T_6) & 31'sh300; // @[Parameters.scala 137:52]
  assign requestARIO_0_1 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_10 = auto_in_ar_bits_addr ^ 30'h200; // @[Parameters.scala 137:31]
  assign _T_11 = {1'b0,$signed(_T_10)}; // @[Parameters.scala 137:49]
  assign _T_13 = $signed(_T_11) & 31'sh300; // @[Parameters.scala 137:52]
  assign requestARIO_0_2 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_16 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_18 = $signed(_T_16) & 31'sh300; // @[Parameters.scala 137:52]
  assign requestAWIO_0_0 = $signed(_T_18) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_20 = auto_in_aw_bits_addr ^ 30'h100; // @[Parameters.scala 137:31]
  assign _T_21 = {1'b0,$signed(_T_20)}; // @[Parameters.scala 137:49]
  assign _T_23 = $signed(_T_21) & 31'sh300; // @[Parameters.scala 137:52]
  assign requestAWIO_0_1 = $signed(_T_23) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_25 = auto_in_aw_bits_addr ^ 30'h200; // @[Parameters.scala 137:31]
  assign _T_26 = {1'b0,$signed(_T_25)}; // @[Parameters.scala 137:49]
  assign _T_28 = $signed(_T_26) & 31'sh300; // @[Parameters.scala 137:52]
  assign requestAWIO_0_2 = $signed(_T_28) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestROI_0_0 = ~auto_out_0_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_2_0 = ~auto_out_2_r_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_0_0 = ~auto_out_0_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_2_0 = ~auto_out_2_b_bits_id; // @[Parameters.scala 47:9]
  assign _T_30 = {requestAWIO_0_2,requestAWIO_0_1}; // @[Xbar.scala 64:75]
  assign _T_31 = {requestAWIO_0_2,requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  assign requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  assign requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  assign requestWIO_0_2 = awIn_0_io_deq_bits[2]; // @[Xbar.scala 65:73]
  assign _T_39 = {requestARIO_0_2,requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  assign _GEN_22 = {{1'd0}, _T_39[2]}; // @[OneHot.scala 32:28]
  assign _T_43 = _GEN_22 | _T_39[1:0]; // @[OneHot.scala 32:28]
  assign _T_45 = {_T_39[2],_T_43[1]}; // @[Cat.scala 29:58]
  assign _GEN_23 = {{1'd0}, _T_31[2]}; // @[OneHot.scala 32:28]
  assign _T_51 = _GEN_23 | _T_31[1:0]; // @[OneHot.scala 32:28]
  assign _T_53 = {_T_31[2],_T_51[1]}; // @[Cat.scala 29:58]
  assign _T_132 = requestARIO_0_0 & auto_out_0_ar_ready; // @[Mux.scala 27:72]
  assign _T_133 = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  assign _T_135 = _T_132 | _T_133; // @[Mux.scala 27:72]
  assign _T_134 = requestARIO_0_2 & auto_out_2_ar_ready; // @[Mux.scala 27:72]
  assign in_0_ar_ready = _T_135 | _T_134; // @[Mux.scala 27:72]
  assign _T_78 = _T_59 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_77 = _T_60 == _T_45; // @[Xbar.scala 111:75]
  assign _T_79 = _T_78 | _T_77; // @[Xbar.scala 112:34]
  assign _T_80 = _T_59 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_82 = _T_79 & _T_80; // @[Xbar.scala 112:48]
  assign io_in_0_ar_ready = in_0_ar_ready & _T_82; // @[Xbar.scala 130:45]
  assign _T_54 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  assign _T_159 = auto_out_0_r_valid & requestROI_0_0; // @[Xbar.scala 222:40]
  assign _T_161 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  assign _T_303 = _T_159 | _T_161; // @[Xbar.scala 246:36]
  assign _T_163 = auto_out_2_r_valid & requestROI_2_0; // @[Xbar.scala 222:40]
  assign _T_304 = _T_303 | _T_163; // @[Xbar.scala 246:36]
  assign _T_380 = _T_373_0 & _T_159; // @[Mux.scala 27:72]
  assign _T_381 = _T_373_1 & _T_161; // @[Mux.scala 27:72]
  assign _T_383 = _T_380 | _T_381; // @[Mux.scala 27:72]
  assign _T_382 = _T_373_2 & _T_163; // @[Mux.scala 27:72]
  assign _T_384 = _T_383 | _T_382; // @[Mux.scala 27:72]
  assign in_0_r_valid = _T_302 ? _T_304 : _T_384; // @[Xbar.scala 278:22]
  assign _T_56 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  assign _T_306 = {_T_163,_T_161,_T_159}; // @[Cat.scala 29:58]
  assign _T_314 = ~_T_313; // @[Arbiter.scala 21:30]
  assign _T_315 = _T_306 & _T_314; // @[Arbiter.scala 21:28]
  assign _T_316 = {_T_315,_T_163,_T_161,_T_159}; // @[Cat.scala 29:58]
  assign _GEN_24 = {{1'd0}, _T_316[5:1]}; // @[package.scala 208:43]
  assign _T_318 = _T_316 | _GEN_24; // @[package.scala 208:43]
  assign _GEN_25 = {{2'd0}, _T_318[5:2]}; // @[package.scala 208:43]
  assign _T_320 = _T_318 | _GEN_25; // @[package.scala 208:43]
  assign _T_323 = {_T_313, 3'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_26 = {{1'd0}, _T_320[5:1]}; // @[Arbiter.scala 22:58]
  assign _T_324 = _GEN_26 | _T_323; // @[Arbiter.scala 22:58]
  assign _T_327 = _T_324[5:3] & _T_324[2:0]; // @[Arbiter.scala 23:39]
  assign _T_328 = ~_T_327; // @[Arbiter.scala 23:18]
  assign _T_344 = _T_328[0] & _T_159; // @[Xbar.scala 250:63]
  assign _T_374_0 = _T_302 ? _T_344 : _T_373_0; // @[Xbar.scala 262:23]
  assign _T_389 = {auto_out_0_r_bits_id,auto_out_0_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  assign _T_390 = _T_374_0 ? _T_389 : 36'h0; // @[Mux.scala 27:72]
  assign _T_345 = _T_328[1] & _T_161; // @[Xbar.scala 250:63]
  assign _T_374_1 = _T_302 ? _T_345 : _T_373_1; // @[Xbar.scala 262:23]
  assign _T_393 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  assign _T_394 = _T_374_1 ? _T_393 : 36'h0; // @[Mux.scala 27:72]
  assign _T_399 = _T_390 | _T_394; // @[Mux.scala 27:72]
  assign _T_346 = _T_328[2] & _T_163; // @[Xbar.scala 250:63]
  assign _T_374_2 = _T_302 ? _T_346 : _T_373_2; // @[Xbar.scala 262:23]
  assign _T_397 = {auto_out_2_r_bits_id,auto_out_2_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  assign _T_398 = _T_374_2 ? _T_397 : 36'h0; // @[Mux.scala 27:72]
  assign _T_400 = _T_399 | _T_398; // @[Mux.scala 27:72]
  assign in_0_r_bits_last = _T_400[0]; // @[Mux.scala 27:72]
  assign _T_58 = _T_56 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  assign _GEN_27 = {{2'd0}, _T_54}; // @[Xbar.scala 106:30]
  assign _T_62 = _T_59 + _GEN_27; // @[Xbar.scala 106:30]
  assign _GEN_28 = {{2'd0}, _T_58}; // @[Xbar.scala 106:48]
  assign _T_64 = _T_62 - _GEN_28; // @[Xbar.scala 106:48]
  assign _T_65 = ~_T_58; // @[Xbar.scala 107:23]
  assign _T_66 = _T_59 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_67 = _T_65 | _T_66; // @[Xbar.scala 107:34]
  assign _T_69 = _T_67 | reset; // @[Xbar.scala 107:22]
  assign _T_70 = ~_T_69; // @[Xbar.scala 107:22]
  assign _T_71 = ~_T_54; // @[Xbar.scala 108:23]
  assign _T_73 = _T_71 | _T_80; // @[Xbar.scala 108:34]
  assign _T_75 = _T_73 | reset; // @[Xbar.scala 108:22]
  assign _T_76 = ~_T_75; // @[Xbar.scala 108:22]
  assign _T_142 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  assign _T_143 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  assign _T_145 = _T_142 | _T_143; // @[Mux.scala 27:72]
  assign _T_144 = requestAWIO_0_2 & auto_out_2_aw_ready; // @[Mux.scala 27:72]
  assign in_0_aw_ready = _T_145 | _T_144; // @[Mux.scala 27:72]
  assign _T_117 = _T_113 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  assign _T_118 = in_0_aw_ready & _T_117; // @[Xbar.scala 139:45]
  assign _T_106 = _T_87 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_105 = _T_88 == _T_53; // @[Xbar.scala 111:75]
  assign _T_107 = _T_106 | _T_105; // @[Xbar.scala 112:34]
  assign _T_108 = _T_87 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_110 = _T_107 & _T_108; // @[Xbar.scala 112:48]
  assign io_in_0_aw_ready = _T_118 & _T_110; // @[Xbar.scala 139:82]
  assign _T_83 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  assign _T_165 = auto_out_0_b_valid & requestBOI_0_0; // @[Xbar.scala 222:40]
  assign _T_167 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  assign _T_408 = _T_165 | _T_167; // @[Xbar.scala 246:36]
  assign _T_169 = auto_out_2_b_valid & requestBOI_2_0; // @[Xbar.scala 222:40]
  assign _T_409 = _T_408 | _T_169; // @[Xbar.scala 246:36]
  assign _T_485 = _T_478_0 & _T_165; // @[Mux.scala 27:72]
  assign _T_486 = _T_478_1 & _T_167; // @[Mux.scala 27:72]
  assign _T_488 = _T_485 | _T_486; // @[Mux.scala 27:72]
  assign _T_487 = _T_478_2 & _T_169; // @[Mux.scala 27:72]
  assign _T_489 = _T_488 | _T_487; // @[Mux.scala 27:72]
  assign in_0_b_valid = _T_407 ? _T_409 : _T_489; // @[Xbar.scala 278:22]
  assign _T_85 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = {{2'd0}, _T_83}; // @[Xbar.scala 106:30]
  assign _T_90 = _T_87 + _GEN_29; // @[Xbar.scala 106:30]
  assign _GEN_30 = {{2'd0}, _T_85}; // @[Xbar.scala 106:48]
  assign _T_92 = _T_90 - _GEN_30; // @[Xbar.scala 106:48]
  assign _T_93 = ~_T_85; // @[Xbar.scala 107:23]
  assign _T_94 = _T_87 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_95 = _T_93 | _T_94; // @[Xbar.scala 107:34]
  assign _T_97 = _T_95 | reset; // @[Xbar.scala 107:22]
  assign _T_98 = ~_T_97; // @[Xbar.scala 107:22]
  assign _T_99 = ~_T_83; // @[Xbar.scala 108:23]
  assign _T_101 = _T_99 | _T_108; // @[Xbar.scala 108:34]
  assign _T_103 = _T_101 | reset; // @[Xbar.scala 108:22]
  assign _T_104 = ~_T_103; // @[Xbar.scala 108:22]
  assign in_0_ar_valid = auto_in_ar_valid & _T_82; // @[Xbar.scala 129:45]
  assign _T_115 = auto_in_aw_valid & _T_117; // @[Xbar.scala 138:45]
  assign in_0_aw_valid = _T_115 & _T_110; // @[Xbar.scala 138:82]
  assign _T_120 = ~_T_113; // @[Xbar.scala 140:54]
  assign _T_122 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_122 | _T_113; // @[Xbar.scala 141:38]
  assign _T_123 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  assign in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  assign _T_152 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  assign _T_153 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  assign _T_155 = _T_152 | _T_153; // @[Mux.scala 27:72]
  assign _T_154 = requestWIO_0_2 & auto_out_2_w_ready; // @[Mux.scala 27:72]
  assign in_0_w_ready = _T_155 | _T_154; // @[Mux.scala 27:72]
  assign _T_126 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  assign out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  assign out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[Xbar.scala 222:40]
  assign out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  assign out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[Xbar.scala 222:40]
  assign _T_176 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  assign _T_182 = _T_176 | out_0_aw_valid; // @[Xbar.scala 258:23]
  assign _T_184 = _T_182 | reset; // @[Xbar.scala 258:12]
  assign _T_185 = ~_T_184; // @[Xbar.scala 258:12]
  assign _T_197 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  assign _T_203 = _T_197 | out_0_ar_valid; // @[Xbar.scala 258:23]
  assign _T_205 = _T_203 | reset; // @[Xbar.scala 258:12]
  assign _T_206 = ~_T_205; // @[Xbar.scala 258:12]
  assign _T_220 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  assign _T_226 = _T_220 | out_1_aw_valid; // @[Xbar.scala 258:23]
  assign _T_228 = _T_226 | reset; // @[Xbar.scala 258:12]
  assign _T_229 = ~_T_228; // @[Xbar.scala 258:12]
  assign _T_241 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  assign _T_247 = _T_241 | out_1_ar_valid; // @[Xbar.scala 258:23]
  assign _T_249 = _T_247 | reset; // @[Xbar.scala 258:12]
  assign _T_250 = ~_T_249; // @[Xbar.scala 258:12]
  assign _T_264 = ~out_2_aw_valid; // @[Xbar.scala 256:60]
  assign _T_270 = _T_264 | out_2_aw_valid; // @[Xbar.scala 258:23]
  assign _T_272 = _T_270 | reset; // @[Xbar.scala 258:12]
  assign _T_273 = ~_T_272; // @[Xbar.scala 258:12]
  assign _T_285 = ~out_2_ar_valid; // @[Xbar.scala 256:60]
  assign _T_291 = _T_285 | out_2_ar_valid; // @[Xbar.scala 258:23]
  assign _T_293 = _T_291 | reset; // @[Xbar.scala 258:12]
  assign _T_294 = ~_T_293; // @[Xbar.scala 258:12]
  assign _T_329 = _T_306 != 3'h0; // @[Arbiter.scala 24:27]
  assign _T_330 = _T_302 & _T_329; // @[Arbiter.scala 24:18]
  assign _T_331 = _T_328 & _T_306; // @[Arbiter.scala 25:29]
  assign _T_332 = {_T_331, 1'h0}; // @[package.scala 199:48]
  assign _T_334 = _T_331 | _T_332[2:0]; // @[package.scala 199:43]
  assign _T_335 = {_T_334, 2'h0}; // @[package.scala 199:48]
  assign _T_337 = _T_334 | _T_335[2:0]; // @[package.scala 199:43]
  assign _T_349 = _T_344 | _T_345; // @[Xbar.scala 255:50]
  assign _T_350 = _T_349 | _T_346; // @[Xbar.scala 255:50]
  assign _T_352 = ~_T_344; // @[Xbar.scala 256:60]
  assign _T_355 = ~_T_345; // @[Xbar.scala 256:60]
  assign _T_356 = _T_352 | _T_355; // @[Xbar.scala 256:57]
  assign _T_357 = ~_T_349; // @[Xbar.scala 256:54]
  assign _T_358 = ~_T_346; // @[Xbar.scala 256:60]
  assign _T_359 = _T_357 | _T_358; // @[Xbar.scala 256:57]
  assign _T_361 = _T_356 & _T_359; // @[Xbar.scala 256:75]
  assign _T_363 = _T_361 | reset; // @[Xbar.scala 256:11]
  assign _T_364 = ~_T_363; // @[Xbar.scala 256:11]
  assign _T_365 = ~_T_304; // @[Xbar.scala 258:13]
  assign _T_368 = _T_365 | _T_350; // @[Xbar.scala 258:23]
  assign _T_370 = _T_368 | reset; // @[Xbar.scala 258:12]
  assign _T_371 = ~_T_370; // @[Xbar.scala 258:12]
  assign _GEN_17 = _T_304 ? 1'h0 : _T_302; // @[Xbar.scala 266:21]
  assign _GEN_18 = _T_56 | _GEN_17; // @[Xbar.scala 267:24]
  assign _T_376_0 = _T_302 ? _T_328[0] : _T_373_0; // @[Xbar.scala 270:24]
  assign _T_376_1 = _T_302 ? _T_328[1] : _T_373_1; // @[Xbar.scala 270:24]
  assign _T_376_2 = _T_302 ? _T_328[2] : _T_373_2; // @[Xbar.scala 270:24]
  assign _T_411 = {_T_169,_T_167,_T_165}; // @[Cat.scala 29:58]
  assign _T_419 = ~_T_418; // @[Arbiter.scala 21:30]
  assign _T_420 = _T_411 & _T_419; // @[Arbiter.scala 21:28]
  assign _T_421 = {_T_420,_T_169,_T_167,_T_165}; // @[Cat.scala 29:58]
  assign _GEN_31 = {{1'd0}, _T_421[5:1]}; // @[package.scala 208:43]
  assign _T_423 = _T_421 | _GEN_31; // @[package.scala 208:43]
  assign _GEN_32 = {{2'd0}, _T_423[5:2]}; // @[package.scala 208:43]
  assign _T_425 = _T_423 | _GEN_32; // @[package.scala 208:43]
  assign _T_428 = {_T_418, 3'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_33 = {{1'd0}, _T_425[5:1]}; // @[Arbiter.scala 22:58]
  assign _T_429 = _GEN_33 | _T_428; // @[Arbiter.scala 22:58]
  assign _T_432 = _T_429[5:3] & _T_429[2:0]; // @[Arbiter.scala 23:39]
  assign _T_433 = ~_T_432; // @[Arbiter.scala 23:18]
  assign _T_434 = _T_411 != 3'h0; // @[Arbiter.scala 24:27]
  assign _T_435 = _T_407 & _T_434; // @[Arbiter.scala 24:18]
  assign _T_436 = _T_433 & _T_411; // @[Arbiter.scala 25:29]
  assign _T_437 = {_T_436, 1'h0}; // @[package.scala 199:48]
  assign _T_439 = _T_436 | _T_437[2:0]; // @[package.scala 199:43]
  assign _T_440 = {_T_439, 2'h0}; // @[package.scala 199:48]
  assign _T_442 = _T_439 | _T_440[2:0]; // @[package.scala 199:43]
  assign _T_449 = _T_433[0] & _T_165; // @[Xbar.scala 250:63]
  assign _T_450 = _T_433[1] & _T_167; // @[Xbar.scala 250:63]
  assign _T_451 = _T_433[2] & _T_169; // @[Xbar.scala 250:63]
  assign _T_454 = _T_449 | _T_450; // @[Xbar.scala 255:50]
  assign _T_455 = _T_454 | _T_451; // @[Xbar.scala 255:50]
  assign _T_457 = ~_T_449; // @[Xbar.scala 256:60]
  assign _T_460 = ~_T_450; // @[Xbar.scala 256:60]
  assign _T_461 = _T_457 | _T_460; // @[Xbar.scala 256:57]
  assign _T_462 = ~_T_454; // @[Xbar.scala 256:54]
  assign _T_463 = ~_T_451; // @[Xbar.scala 256:60]
  assign _T_464 = _T_462 | _T_463; // @[Xbar.scala 256:57]
  assign _T_466 = _T_461 & _T_464; // @[Xbar.scala 256:75]
  assign _T_468 = _T_466 | reset; // @[Xbar.scala 256:11]
  assign _T_469 = ~_T_468; // @[Xbar.scala 256:11]
  assign _T_470 = ~_T_409; // @[Xbar.scala 258:13]
  assign _T_473 = _T_470 | _T_455; // @[Xbar.scala 258:23]
  assign _T_475 = _T_473 | reset; // @[Xbar.scala 258:12]
  assign _T_476 = ~_T_475; // @[Xbar.scala 258:12]
  assign _T_479_0 = _T_407 ? _T_449 : _T_478_0; // @[Xbar.scala 262:23]
  assign _T_479_1 = _T_407 ? _T_450 : _T_478_1; // @[Xbar.scala 262:23]
  assign _T_479_2 = _T_407 ? _T_451 : _T_478_2; // @[Xbar.scala 262:23]
  assign _GEN_20 = _T_409 ? 1'h0 : _T_407; // @[Xbar.scala 266:21]
  assign _GEN_21 = _T_85 | _GEN_20; // @[Xbar.scala 267:24]
  assign _T_481_0 = _T_407 ? _T_433[0] : _T_478_0; // @[Xbar.scala 270:24]
  assign _T_481_1 = _T_407 ? _T_433[1] : _T_478_1; // @[Xbar.scala 270:24]
  assign _T_481_2 = _T_407 ? _T_433[2] : _T_478_2; // @[Xbar.scala 270:24]
  assign _T_492 = {auto_out_0_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  assign _T_493 = _T_479_0 ? _T_492 : 3'h0; // @[Mux.scala 27:72]
  assign _T_494 = {auto_out_1_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  assign _T_495 = _T_479_1 ? _T_494 : 3'h0; // @[Mux.scala 27:72]
  assign _T_496 = {auto_out_2_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  assign _T_497 = _T_479_2 ? _T_496 : 3'h0; // @[Mux.scala 27:72]
  assign _T_498 = _T_493 | _T_495; // @[Mux.scala 27:72]
  assign _T_499 = _T_498 | _T_497; // @[Mux.scala 27:72]
  assign auto_in_aw_ready = _T_118 & _T_110; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_407 ? _T_409 : _T_489; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_499[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_82; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_302 ? _T_304 : _T_384; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_400[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_400[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_400[0]; // @[LazyModule.scala 173:31]
  assign auto_out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_valid = in_0_w_valid & requestWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_2_b_ready = auto_in_b_ready & _T_481_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_2_r_ready = auto_in_r_ready & _T_376_2; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_481_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_376_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_481_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_r_ready = auto_in_r_ready & _T_376_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_120; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {_T_30,requestAWIO_0_0}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_126 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_59 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_60 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_302 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_373_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_373_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_373_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_313 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_113 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_87 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_88 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_407 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_478_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_478_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_478_2 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_418 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_59 <= 3'h0;
    end else begin
      _T_59 <= _T_64;
    end
    if (_T_54) begin
      _T_60 <= _T_45;
    end
    _T_302 <= reset | _GEN_18;
    if (reset) begin
      _T_373_0 <= 1'h0;
    end else if (_T_302) begin
      _T_373_0 <= _T_344;
    end
    if (reset) begin
      _T_373_1 <= 1'h0;
    end else if (_T_302) begin
      _T_373_1 <= _T_345;
    end
    if (reset) begin
      _T_373_2 <= 1'h0;
    end else if (_T_302) begin
      _T_373_2 <= _T_346;
    end
    if (reset) begin
      _T_313 <= 3'h7;
    end else if (_T_330) begin
      _T_313 <= _T_337;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else if (_T_123) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _GEN_2;
    end
    if (reset) begin
      _T_87 <= 3'h0;
    end else begin
      _T_87 <= _T_92;
    end
    if (_T_83) begin
      _T_88 <= _T_53;
    end
    _T_407 <= reset | _GEN_21;
    if (reset) begin
      _T_478_0 <= 1'h0;
    end else if (_T_407) begin
      _T_478_0 <= _T_449;
    end
    if (reset) begin
      _T_478_1 <= 1'h0;
    end else if (_T_407) begin
      _T_478_1 <= _T_450;
    end
    if (reset) begin
      _T_478_2 <= 1'h0;
    end else if (_T_407) begin
      _T_478_2 <= _T_451;
    end
    if (reset) begin
      _T_418 <= 3'h7;
    end else if (_T_435) begin
      _T_418 <= _T_442;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_70) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_70) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_76) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_76) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_98) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_104) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_185) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_185) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_206) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_206) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_229) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_229) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_250) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_250) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_273) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_273) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_294) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_294) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_364) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_364) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_371) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_371) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_469) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_469) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_476) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_476) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BundleBridgeToAXI4(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49]
endmodule
module AXI4StreamToBundleBridge(
  output        auto_in_ready,
  input         auto_in_valid,
  input  [15:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [15:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module BundleBridgeToAXI4Stream(
  output       auto_in_ready,
  input        auto_in_valid,
  input  [7:0] auto_in_bits_data,
  input        auto_in_bits_last,
  input        auto_out_ready,
  output       auto_out_valid,
  output [7:0] auto_out_bits_data,
  output       auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module AXI4HyperSpace(
  input         clock,
  input         reset,
  output        ioMem_0_aw_ready,
  input         ioMem_0_aw_valid,
  input         ioMem_0_aw_bits_id,
  input  [31:0] ioMem_0_aw_bits_addr,
  input  [7:0]  ioMem_0_aw_bits_len,
  input  [2:0]  ioMem_0_aw_bits_size,
  input  [1:0]  ioMem_0_aw_bits_burst,
  input         ioMem_0_aw_bits_lock,
  input  [3:0]  ioMem_0_aw_bits_cache,
  input  [2:0]  ioMem_0_aw_bits_prot,
  input  [3:0]  ioMem_0_aw_bits_qos,
  output        ioMem_0_w_ready,
  input         ioMem_0_w_valid,
  input  [31:0] ioMem_0_w_bits_data,
  input  [3:0]  ioMem_0_w_bits_strb,
  input         ioMem_0_w_bits_last,
  input         ioMem_0_b_ready,
  output        ioMem_0_b_valid,
  output        ioMem_0_b_bits_id,
  output [1:0]  ioMem_0_b_bits_resp,
  output        ioMem_0_ar_ready,
  input         ioMem_0_ar_valid,
  input         ioMem_0_ar_bits_id,
  input  [31:0] ioMem_0_ar_bits_addr,
  input  [7:0]  ioMem_0_ar_bits_len,
  input  [2:0]  ioMem_0_ar_bits_size,
  input  [1:0]  ioMem_0_ar_bits_burst,
  input         ioMem_0_ar_bits_lock,
  input  [3:0]  ioMem_0_ar_bits_cache,
  input  [2:0]  ioMem_0_ar_bits_prot,
  input  [3:0]  ioMem_0_ar_bits_qos,
  input         ioMem_0_r_ready,
  output        ioMem_0_r_valid,
  output        ioMem_0_r_bits_id,
  output [31:0] ioMem_0_r_bits_data,
  output [1:0]  ioMem_0_r_bits_resp,
  output        ioMem_0_r_bits_last,
  output        in_0_ready,
  input         in_0_valid,
  input  [7:0]  in_0_bits_data,
  input         in_0_bits_last,
  input         out_0_ready,
  output        out_0_valid,
  output [15:0] out_0_bits_data,
  output        out_0_bits_last
);
  wire  widthAdapter_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  fft_clock; // @[HyperSpace.scala 62:76]
  wire  fft_reset; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_aw_ready; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_aw_valid; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_aw_bits_id; // @[HyperSpace.scala 62:76]
  wire [29:0] fft_auto_mem_in_aw_bits_addr; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_w_ready; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_w_valid; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_b_ready; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_b_valid; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_b_bits_id; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_ar_ready; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_ar_valid; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_ar_bits_id; // @[HyperSpace.scala 62:76]
  wire [29:0] fft_auto_mem_in_ar_bits_addr; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_r_ready; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_r_valid; // @[HyperSpace.scala 62:76]
  wire  fft_auto_mem_in_r_bits_id; // @[HyperSpace.scala 62:76]
  wire [31:0] fft_auto_mem_in_r_bits_data; // @[HyperSpace.scala 62:76]
  wire  fft_auto_stream_in_ready; // @[HyperSpace.scala 62:76]
  wire  fft_auto_stream_in_valid; // @[HyperSpace.scala 62:76]
  wire [31:0] fft_auto_stream_in_bits_data; // @[HyperSpace.scala 62:76]
  wire  fft_auto_stream_in_bits_last; // @[HyperSpace.scala 62:76]
  wire  fft_auto_stream_out_ready; // @[HyperSpace.scala 62:76]
  wire  fft_auto_stream_out_valid; // @[HyperSpace.scala 62:76]
  wire [31:0] fft_auto_stream_out_bits_data; // @[HyperSpace.scala 62:76]
  wire  fft_auto_stream_out_bits_last; // @[HyperSpace.scala 62:76]
  wire  mag_clock; // @[HyperSpace.scala 63:76]
  wire  mag_reset; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_aw_ready; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_aw_valid; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_aw_bits_id; // @[HyperSpace.scala 63:76]
  wire [29:0] mag_auto_mem_in_aw_bits_addr; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_w_ready; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_w_valid; // @[HyperSpace.scala 63:76]
  wire [31:0] mag_auto_mem_in_w_bits_data; // @[HyperSpace.scala 63:76]
  wire [3:0] mag_auto_mem_in_w_bits_strb; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_b_ready; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_b_valid; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_b_bits_id; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_ar_ready; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_ar_valid; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_ar_bits_id; // @[HyperSpace.scala 63:76]
  wire [29:0] mag_auto_mem_in_ar_bits_addr; // @[HyperSpace.scala 63:76]
  wire [2:0] mag_auto_mem_in_ar_bits_size; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_r_ready; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_r_valid; // @[HyperSpace.scala 63:76]
  wire  mag_auto_mem_in_r_bits_id; // @[HyperSpace.scala 63:76]
  wire [31:0] mag_auto_mem_in_r_bits_data; // @[HyperSpace.scala 63:76]
  wire  mag_auto_master_out_ready; // @[HyperSpace.scala 63:76]
  wire  mag_auto_master_out_valid; // @[HyperSpace.scala 63:76]
  wire [15:0] mag_auto_master_out_bits_data; // @[HyperSpace.scala 63:76]
  wire  mag_auto_master_out_bits_last; // @[HyperSpace.scala 63:76]
  wire  mag_auto_slave_in_ready; // @[HyperSpace.scala 63:76]
  wire  mag_auto_slave_in_valid; // @[HyperSpace.scala 63:76]
  wire [31:0] mag_auto_slave_in_bits_data; // @[HyperSpace.scala 63:76]
  wire  mag_auto_slave_in_bits_last; // @[HyperSpace.scala 63:76]
  wire  cfar_clock; // @[HyperSpace.scala 64:76]
  wire  cfar_reset; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_aw_ready; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_aw_valid; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_aw_bits_id; // @[HyperSpace.scala 64:76]
  wire [29:0] cfar_auto_mem_in_aw_bits_addr; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_w_ready; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_w_valid; // @[HyperSpace.scala 64:76]
  wire [31:0] cfar_auto_mem_in_w_bits_data; // @[HyperSpace.scala 64:76]
  wire [3:0] cfar_auto_mem_in_w_bits_strb; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_b_ready; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_b_valid; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_b_bits_id; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_ar_ready; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_ar_valid; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_ar_bits_id; // @[HyperSpace.scala 64:76]
  wire [29:0] cfar_auto_mem_in_ar_bits_addr; // @[HyperSpace.scala 64:76]
  wire [2:0] cfar_auto_mem_in_ar_bits_size; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_r_ready; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_r_valid; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_mem_in_r_bits_id; // @[HyperSpace.scala 64:76]
  wire [31:0] cfar_auto_mem_in_r_bits_data; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_master_out_ready; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_master_out_valid; // @[HyperSpace.scala 64:76]
  wire [47:0] cfar_auto_master_out_bits_data; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_master_out_bits_last; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_slave_in_ready; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_slave_in_valid; // @[HyperSpace.scala 64:76]
  wire [15:0] cfar_auto_slave_in_bits_data; // @[HyperSpace.scala 64:76]
  wire  cfar_auto_slave_in_bits_last; // @[HyperSpace.scala 64:76]
  wire  widthAdapter_1_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [47:0] widthAdapter_1_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [15:0] widthAdapter_1_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  buffer_clock; // @[Buffer.scala 29:28]
  wire  buffer_reset; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_clock; // @[Buffer.scala 29:28]
  wire  buffer_1_reset; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_valid; // @[Buffer.scala 29:28]
  wire [15:0] buffer_1_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_valid; // @[Buffer.scala 29:28]
  wire [15:0] buffer_1_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_clock; // @[Buffer.scala 29:28]
  wire  buffer_2_reset; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_clock; // @[Buffer.scala 29:28]
  wire  buffer_3_reset; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_valid; // @[Buffer.scala 29:28]
  wire [47:0] buffer_3_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_valid; // @[Buffer.scala 29:28]
  wire [47:0] buffer_3_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  bus_clock; // @[HyperSpace.scala 49:58]
  wire  bus_reset; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_aw_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_aw_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_aw_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_in_aw_bits_addr; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_w_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_w_valid; // @[HyperSpace.scala 49:58]
  wire [31:0] bus_auto_in_w_bits_data; // @[HyperSpace.scala 49:58]
  wire [3:0] bus_auto_in_w_bits_strb; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_w_bits_last; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_b_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_b_valid; // @[HyperSpace.scala 49:58]
  wire [1:0] bus_auto_in_b_bits_resp; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_ar_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_ar_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_ar_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_in_ar_bits_addr; // @[HyperSpace.scala 49:58]
  wire [2:0] bus_auto_in_ar_bits_size; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_r_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_r_valid; // @[HyperSpace.scala 49:58]
  wire [31:0] bus_auto_in_r_bits_data; // @[HyperSpace.scala 49:58]
  wire [1:0] bus_auto_in_r_bits_resp; // @[HyperSpace.scala 49:58]
  wire  bus_auto_in_r_bits_last; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_aw_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_aw_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_aw_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_out_2_aw_bits_addr; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_w_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_w_valid; // @[HyperSpace.scala 49:58]
  wire [31:0] bus_auto_out_2_w_bits_data; // @[HyperSpace.scala 49:58]
  wire [3:0] bus_auto_out_2_w_bits_strb; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_b_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_b_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_b_bits_id; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_ar_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_ar_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_ar_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_out_2_ar_bits_addr; // @[HyperSpace.scala 49:58]
  wire [2:0] bus_auto_out_2_ar_bits_size; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_r_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_r_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_2_r_bits_id; // @[HyperSpace.scala 49:58]
  wire [31:0] bus_auto_out_2_r_bits_data; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_aw_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_aw_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_aw_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_out_1_aw_bits_addr; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_w_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_w_valid; // @[HyperSpace.scala 49:58]
  wire [31:0] bus_auto_out_1_w_bits_data; // @[HyperSpace.scala 49:58]
  wire [3:0] bus_auto_out_1_w_bits_strb; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_b_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_b_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_b_bits_id; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_ar_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_ar_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_ar_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_out_1_ar_bits_addr; // @[HyperSpace.scala 49:58]
  wire [2:0] bus_auto_out_1_ar_bits_size; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_r_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_r_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_1_r_bits_id; // @[HyperSpace.scala 49:58]
  wire [31:0] bus_auto_out_1_r_bits_data; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_aw_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_aw_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_aw_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_out_0_aw_bits_addr; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_w_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_w_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_b_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_b_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_b_bits_id; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_ar_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_ar_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_ar_bits_id; // @[HyperSpace.scala 49:58]
  wire [29:0] bus_auto_out_0_ar_bits_addr; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_r_ready; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_r_valid; // @[HyperSpace.scala 49:58]
  wire  bus_auto_out_0_r_bits_id; // @[HyperSpace.scala 49:58]
  wire [31:0] bus_auto_out_0_r_bits_data; // @[HyperSpace.scala 49:58]
  wire  converter_auto_in_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_aw_bits_addr; // @[Node.scala 65:31]
  wire  converter_auto_in_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_in_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_in_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_in_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_in_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_in_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_r_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_aw_bits_addr; // @[Node.scala 65:31]
  wire  converter_auto_out_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_out_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_out_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_out_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_out_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_r_bits_last; // @[Node.scala 65:31]
  wire  converter_1_auto_in_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_valid; // @[Nodes.scala 165:31]
  wire [15:0] converter_1_auto_in_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_bits_last; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_valid; // @[Nodes.scala 165:31]
  wire [15:0] converter_1_auto_out_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_bits_last; // @[Nodes.scala 165:31]
  wire  converter_2_auto_in_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_in_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_bits_last; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_out_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_bits_last; // @[Nodes.scala 201:31]
  AXI4StreamWidthAdapater_4_to_1 widthAdapter ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_clock),
    .reset(widthAdapter_reset),
    .auto_in_ready(widthAdapter_auto_in_ready),
    .auto_in_valid(widthAdapter_auto_in_valid),
    .auto_in_bits_data(widthAdapter_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_auto_in_bits_last),
    .auto_out_ready(widthAdapter_auto_out_ready),
    .auto_out_valid(widthAdapter_auto_out_valid),
    .auto_out_bits_data(widthAdapter_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_auto_out_bits_last)
  );
  AXI4FFTBlock fft ( // @[HyperSpace.scala 62:76]
    .clock(fft_clock),
    .reset(fft_reset),
    .auto_mem_in_aw_ready(fft_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(fft_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(fft_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(fft_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(fft_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(fft_auto_mem_in_w_valid),
    .auto_mem_in_b_ready(fft_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(fft_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(fft_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(fft_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(fft_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(fft_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(fft_auto_mem_in_ar_bits_addr),
    .auto_mem_in_r_ready(fft_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(fft_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(fft_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(fft_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(fft_auto_stream_in_ready),
    .auto_stream_in_valid(fft_auto_stream_in_valid),
    .auto_stream_in_bits_data(fft_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(fft_auto_stream_in_bits_last),
    .auto_stream_out_ready(fft_auto_stream_out_ready),
    .auto_stream_out_valid(fft_auto_stream_out_valid),
    .auto_stream_out_bits_data(fft_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(fft_auto_stream_out_bits_last)
  );
  AXI4LogMagMuxBlock mag ( // @[HyperSpace.scala 63:76]
    .clock(mag_clock),
    .reset(mag_reset),
    .auto_mem_in_aw_ready(mag_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(mag_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(mag_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(mag_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(mag_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(mag_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(mag_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(mag_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(mag_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(mag_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(mag_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(mag_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(mag_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(mag_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(mag_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(mag_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(mag_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(mag_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(mag_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(mag_auto_mem_in_r_bits_data),
    .auto_master_out_ready(mag_auto_master_out_ready),
    .auto_master_out_valid(mag_auto_master_out_valid),
    .auto_master_out_bits_data(mag_auto_master_out_bits_data),
    .auto_master_out_bits_last(mag_auto_master_out_bits_last),
    .auto_slave_in_ready(mag_auto_slave_in_ready),
    .auto_slave_in_valid(mag_auto_slave_in_valid),
    .auto_slave_in_bits_data(mag_auto_slave_in_bits_data),
    .auto_slave_in_bits_last(mag_auto_slave_in_bits_last)
  );
  AXI4CFARBlock cfar ( // @[HyperSpace.scala 64:76]
    .clock(cfar_clock),
    .reset(cfar_reset),
    .auto_mem_in_aw_ready(cfar_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(cfar_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(cfar_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(cfar_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(cfar_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(cfar_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(cfar_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(cfar_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(cfar_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(cfar_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(cfar_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(cfar_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(cfar_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(cfar_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(cfar_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(cfar_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(cfar_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(cfar_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(cfar_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(cfar_auto_mem_in_r_bits_data),
    .auto_master_out_ready(cfar_auto_master_out_ready),
    .auto_master_out_valid(cfar_auto_master_out_valid),
    .auto_master_out_bits_data(cfar_auto_master_out_bits_data),
    .auto_master_out_bits_last(cfar_auto_master_out_bits_last),
    .auto_slave_in_ready(cfar_auto_slave_in_ready),
    .auto_slave_in_valid(cfar_auto_slave_in_valid),
    .auto_slave_in_bits_data(cfar_auto_slave_in_bits_data),
    .auto_slave_in_bits_last(cfar_auto_slave_in_bits_last)
  );
  AXI4StreamWidthAdapater_1_to_3 widthAdapter_1 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_1_clock),
    .reset(widthAdapter_1_reset),
    .auto_in_ready(widthAdapter_1_auto_in_ready),
    .auto_in_valid(widthAdapter_1_auto_in_valid),
    .auto_in_bits_data(widthAdapter_1_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_1_auto_in_bits_last),
    .auto_out_ready(widthAdapter_1_auto_out_ready),
    .auto_out_valid(widthAdapter_1_auto_out_valid),
    .auto_out_bits_data(widthAdapter_1_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_1_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer ( // @[Buffer.scala 29:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_ready(buffer_auto_in_ready),
    .auto_in_valid(buffer_auto_in_valid),
    .auto_in_bits_data(buffer_auto_in_bits_data),
    .auto_in_bits_last(buffer_auto_in_bits_last),
    .auto_out_ready(buffer_auto_out_ready),
    .auto_out_valid(buffer_auto_out_valid),
    .auto_out_bits_data(buffer_auto_out_bits_data),
    .auto_out_bits_last(buffer_auto_out_bits_last)
  );
  AXI4StreamBuffer_1 buffer_1 ( // @[Buffer.scala 29:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_ready(buffer_1_auto_in_ready),
    .auto_in_valid(buffer_1_auto_in_valid),
    .auto_in_bits_data(buffer_1_auto_in_bits_data),
    .auto_in_bits_last(buffer_1_auto_in_bits_last),
    .auto_out_ready(buffer_1_auto_out_ready),
    .auto_out_valid(buffer_1_auto_out_valid),
    .auto_out_bits_data(buffer_1_auto_out_bits_data),
    .auto_out_bits_last(buffer_1_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_2 ( // @[Buffer.scala 29:28]
    .clock(buffer_2_clock),
    .reset(buffer_2_reset),
    .auto_in_ready(buffer_2_auto_in_ready),
    .auto_in_valid(buffer_2_auto_in_valid),
    .auto_in_bits_data(buffer_2_auto_in_bits_data),
    .auto_in_bits_last(buffer_2_auto_in_bits_last),
    .auto_out_ready(buffer_2_auto_out_ready),
    .auto_out_valid(buffer_2_auto_out_valid),
    .auto_out_bits_data(buffer_2_auto_out_bits_data),
    .auto_out_bits_last(buffer_2_auto_out_bits_last)
  );
  AXI4StreamBuffer_3 buffer_3 ( // @[Buffer.scala 29:28]
    .clock(buffer_3_clock),
    .reset(buffer_3_reset),
    .auto_in_ready(buffer_3_auto_in_ready),
    .auto_in_valid(buffer_3_auto_in_valid),
    .auto_in_bits_data(buffer_3_auto_in_bits_data),
    .auto_in_bits_last(buffer_3_auto_in_bits_last),
    .auto_out_ready(buffer_3_auto_out_ready),
    .auto_out_valid(buffer_3_auto_out_valid),
    .auto_out_bits_data(buffer_3_auto_out_bits_data),
    .auto_out_bits_last(buffer_3_auto_out_bits_last)
  );
  AXI4Xbar bus ( // @[HyperSpace.scala 49:58]
    .clock(bus_clock),
    .reset(bus_reset),
    .auto_in_aw_ready(bus_auto_in_aw_ready),
    .auto_in_aw_valid(bus_auto_in_aw_valid),
    .auto_in_aw_bits_id(bus_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(bus_auto_in_aw_bits_addr),
    .auto_in_w_ready(bus_auto_in_w_ready),
    .auto_in_w_valid(bus_auto_in_w_valid),
    .auto_in_w_bits_data(bus_auto_in_w_bits_data),
    .auto_in_w_bits_strb(bus_auto_in_w_bits_strb),
    .auto_in_w_bits_last(bus_auto_in_w_bits_last),
    .auto_in_b_ready(bus_auto_in_b_ready),
    .auto_in_b_valid(bus_auto_in_b_valid),
    .auto_in_b_bits_resp(bus_auto_in_b_bits_resp),
    .auto_in_ar_ready(bus_auto_in_ar_ready),
    .auto_in_ar_valid(bus_auto_in_ar_valid),
    .auto_in_ar_bits_id(bus_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(bus_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(bus_auto_in_ar_bits_size),
    .auto_in_r_ready(bus_auto_in_r_ready),
    .auto_in_r_valid(bus_auto_in_r_valid),
    .auto_in_r_bits_data(bus_auto_in_r_bits_data),
    .auto_in_r_bits_resp(bus_auto_in_r_bits_resp),
    .auto_in_r_bits_last(bus_auto_in_r_bits_last),
    .auto_out_2_aw_ready(bus_auto_out_2_aw_ready),
    .auto_out_2_aw_valid(bus_auto_out_2_aw_valid),
    .auto_out_2_aw_bits_id(bus_auto_out_2_aw_bits_id),
    .auto_out_2_aw_bits_addr(bus_auto_out_2_aw_bits_addr),
    .auto_out_2_w_ready(bus_auto_out_2_w_ready),
    .auto_out_2_w_valid(bus_auto_out_2_w_valid),
    .auto_out_2_w_bits_data(bus_auto_out_2_w_bits_data),
    .auto_out_2_w_bits_strb(bus_auto_out_2_w_bits_strb),
    .auto_out_2_b_ready(bus_auto_out_2_b_ready),
    .auto_out_2_b_valid(bus_auto_out_2_b_valid),
    .auto_out_2_b_bits_id(bus_auto_out_2_b_bits_id),
    .auto_out_2_ar_ready(bus_auto_out_2_ar_ready),
    .auto_out_2_ar_valid(bus_auto_out_2_ar_valid),
    .auto_out_2_ar_bits_id(bus_auto_out_2_ar_bits_id),
    .auto_out_2_ar_bits_addr(bus_auto_out_2_ar_bits_addr),
    .auto_out_2_ar_bits_size(bus_auto_out_2_ar_bits_size),
    .auto_out_2_r_ready(bus_auto_out_2_r_ready),
    .auto_out_2_r_valid(bus_auto_out_2_r_valid),
    .auto_out_2_r_bits_id(bus_auto_out_2_r_bits_id),
    .auto_out_2_r_bits_data(bus_auto_out_2_r_bits_data),
    .auto_out_1_aw_ready(bus_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(bus_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(bus_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(bus_auto_out_1_aw_bits_addr),
    .auto_out_1_w_ready(bus_auto_out_1_w_ready),
    .auto_out_1_w_valid(bus_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(bus_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(bus_auto_out_1_w_bits_strb),
    .auto_out_1_b_ready(bus_auto_out_1_b_ready),
    .auto_out_1_b_valid(bus_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(bus_auto_out_1_b_bits_id),
    .auto_out_1_ar_ready(bus_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(bus_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(bus_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(bus_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(bus_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(bus_auto_out_1_r_ready),
    .auto_out_1_r_valid(bus_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(bus_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(bus_auto_out_1_r_bits_data),
    .auto_out_0_aw_ready(bus_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(bus_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_id(bus_auto_out_0_aw_bits_id),
    .auto_out_0_aw_bits_addr(bus_auto_out_0_aw_bits_addr),
    .auto_out_0_w_ready(bus_auto_out_0_w_ready),
    .auto_out_0_w_valid(bus_auto_out_0_w_valid),
    .auto_out_0_b_ready(bus_auto_out_0_b_ready),
    .auto_out_0_b_valid(bus_auto_out_0_b_valid),
    .auto_out_0_b_bits_id(bus_auto_out_0_b_bits_id),
    .auto_out_0_ar_ready(bus_auto_out_0_ar_ready),
    .auto_out_0_ar_valid(bus_auto_out_0_ar_valid),
    .auto_out_0_ar_bits_id(bus_auto_out_0_ar_bits_id),
    .auto_out_0_ar_bits_addr(bus_auto_out_0_ar_bits_addr),
    .auto_out_0_r_ready(bus_auto_out_0_r_ready),
    .auto_out_0_r_valid(bus_auto_out_0_r_valid),
    .auto_out_0_r_bits_id(bus_auto_out_0_r_bits_id),
    .auto_out_0_r_bits_data(bus_auto_out_0_r_bits_data)
  );
  BundleBridgeToAXI4 converter ( // @[Node.scala 65:31]
    .auto_in_aw_ready(converter_auto_in_aw_ready),
    .auto_in_aw_valid(converter_auto_in_aw_valid),
    .auto_in_aw_bits_id(converter_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(converter_auto_in_aw_bits_addr),
    .auto_in_w_ready(converter_auto_in_w_ready),
    .auto_in_w_valid(converter_auto_in_w_valid),
    .auto_in_w_bits_data(converter_auto_in_w_bits_data),
    .auto_in_w_bits_strb(converter_auto_in_w_bits_strb),
    .auto_in_w_bits_last(converter_auto_in_w_bits_last),
    .auto_in_b_ready(converter_auto_in_b_ready),
    .auto_in_b_valid(converter_auto_in_b_valid),
    .auto_in_b_bits_resp(converter_auto_in_b_bits_resp),
    .auto_in_ar_ready(converter_auto_in_ar_ready),
    .auto_in_ar_valid(converter_auto_in_ar_valid),
    .auto_in_ar_bits_id(converter_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(converter_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(converter_auto_in_ar_bits_size),
    .auto_in_r_ready(converter_auto_in_r_ready),
    .auto_in_r_valid(converter_auto_in_r_valid),
    .auto_in_r_bits_data(converter_auto_in_r_bits_data),
    .auto_in_r_bits_resp(converter_auto_in_r_bits_resp),
    .auto_in_r_bits_last(converter_auto_in_r_bits_last),
    .auto_out_aw_ready(converter_auto_out_aw_ready),
    .auto_out_aw_valid(converter_auto_out_aw_valid),
    .auto_out_aw_bits_id(converter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(converter_auto_out_aw_bits_addr),
    .auto_out_w_ready(converter_auto_out_w_ready),
    .auto_out_w_valid(converter_auto_out_w_valid),
    .auto_out_w_bits_data(converter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(converter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(converter_auto_out_w_bits_last),
    .auto_out_b_ready(converter_auto_out_b_ready),
    .auto_out_b_valid(converter_auto_out_b_valid),
    .auto_out_b_bits_resp(converter_auto_out_b_bits_resp),
    .auto_out_ar_ready(converter_auto_out_ar_ready),
    .auto_out_ar_valid(converter_auto_out_ar_valid),
    .auto_out_ar_bits_id(converter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(converter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(converter_auto_out_ar_bits_size),
    .auto_out_r_ready(converter_auto_out_r_ready),
    .auto_out_r_valid(converter_auto_out_r_valid),
    .auto_out_r_bits_data(converter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(converter_auto_out_r_bits_resp),
    .auto_out_r_bits_last(converter_auto_out_r_bits_last)
  );
  AXI4StreamToBundleBridge converter_1 ( // @[Nodes.scala 165:31]
    .auto_in_ready(converter_1_auto_in_ready),
    .auto_in_valid(converter_1_auto_in_valid),
    .auto_in_bits_data(converter_1_auto_in_bits_data),
    .auto_in_bits_last(converter_1_auto_in_bits_last),
    .auto_out_ready(converter_1_auto_out_ready),
    .auto_out_valid(converter_1_auto_out_valid),
    .auto_out_bits_data(converter_1_auto_out_bits_data),
    .auto_out_bits_last(converter_1_auto_out_bits_last)
  );
  BundleBridgeToAXI4Stream converter_2 ( // @[Nodes.scala 201:31]
    .auto_in_ready(converter_2_auto_in_ready),
    .auto_in_valid(converter_2_auto_in_valid),
    .auto_in_bits_data(converter_2_auto_in_bits_data),
    .auto_in_bits_last(converter_2_auto_in_bits_last),
    .auto_out_ready(converter_2_auto_out_ready),
    .auto_out_valid(converter_2_auto_out_valid),
    .auto_out_bits_data(converter_2_auto_out_bits_data),
    .auto_out_bits_last(converter_2_auto_out_bits_last)
  );
  assign ioMem_0_aw_ready = converter_auto_in_aw_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_w_ready = converter_auto_in_w_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_b_valid = converter_auto_in_b_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_resp = converter_auto_in_b_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_ar_ready = converter_auto_in_ar_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_r_valid = converter_auto_in_r_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_data = converter_auto_in_r_bits_data; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_resp = converter_auto_in_r_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_last = converter_auto_in_r_bits_last; // @[Nodes.scala 624:60]
  assign in_0_ready = converter_2_auto_in_ready; // @[Nodes.scala 624:60]
  assign out_0_valid = converter_1_auto_out_valid; // @[Nodes.scala 649:56]
  assign out_0_bits_data = converter_1_auto_out_bits_data; // @[Nodes.scala 649:56]
  assign out_0_bits_last = converter_1_auto_out_bits_last; // @[Nodes.scala 649:56]
  assign widthAdapter_clock = clock;
  assign widthAdapter_reset = reset;
  assign widthAdapter_auto_in_valid = converter_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_data = converter_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_last = converter_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_out_ready = buffer_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_auto_mem_in_aw_valid = bus_auto_out_0_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_id = bus_auto_out_0_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_addr = bus_auto_out_0_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_valid = bus_auto_out_0_w_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_b_ready = bus_auto_out_0_b_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_valid = bus_auto_out_0_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_id = bus_auto_out_0_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_addr = bus_auto_out_0_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_r_ready = bus_auto_out_0_r_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_valid = buffer_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_data = buffer_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_last = buffer_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_out_ready = buffer_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_clock = clock;
  assign mag_reset = reset;
  assign mag_auto_mem_in_aw_valid = bus_auto_out_1_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_id = bus_auto_out_1_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_addr = bus_auto_out_1_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_valid = bus_auto_out_1_w_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_data = bus_auto_out_1_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_strb = bus_auto_out_1_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_b_ready = bus_auto_out_1_b_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_valid = bus_auto_out_1_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_id = bus_auto_out_1_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_addr = bus_auto_out_1_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_size = bus_auto_out_1_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_r_ready = bus_auto_out_1_r_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_master_out_ready = buffer_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_auto_slave_in_valid = buffer_auto_out_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_slave_in_bits_data = buffer_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_slave_in_bits_last = buffer_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign cfar_clock = clock;
  assign cfar_reset = reset;
  assign cfar_auto_mem_in_aw_valid = bus_auto_out_2_aw_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_aw_bits_id = bus_auto_out_2_aw_bits_id; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_aw_bits_addr = bus_auto_out_2_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_w_valid = bus_auto_out_2_w_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_w_bits_data = bus_auto_out_2_w_bits_data; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_w_bits_strb = bus_auto_out_2_w_bits_strb; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_b_ready = bus_auto_out_2_b_ready; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_valid = bus_auto_out_2_ar_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_bits_id = bus_auto_out_2_ar_bits_id; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_bits_addr = bus_auto_out_2_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_ar_bits_size = bus_auto_out_2_ar_bits_size; // @[LazyModule.scala 167:31]
  assign cfar_auto_mem_in_r_ready = bus_auto_out_2_r_ready; // @[LazyModule.scala 167:31]
  assign cfar_auto_master_out_ready = buffer_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign cfar_auto_slave_in_valid = buffer_1_auto_out_valid; // @[LazyModule.scala 167:31]
  assign cfar_auto_slave_in_bits_data = buffer_1_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign cfar_auto_slave_in_bits_last = buffer_1_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_clock = clock;
  assign widthAdapter_1_reset = reset;
  assign widthAdapter_1_auto_in_valid = buffer_3_auto_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_auto_in_bits_data = buffer_3_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_auto_in_bits_last = buffer_3_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_auto_out_ready = converter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_valid = fft_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_data = fft_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_last = fft_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_auto_out_ready = mag_auto_slave_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_1_clock = clock;
  assign buffer_1_reset = reset;
  assign buffer_1_auto_in_valid = mag_auto_master_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_data = mag_auto_master_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_last = mag_auto_master_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_out_ready = cfar_auto_slave_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_2_clock = clock;
  assign buffer_2_reset = reset;
  assign buffer_2_auto_in_valid = widthAdapter_auto_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_data = widthAdapter_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_last = widthAdapter_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_out_ready = fft_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_3_clock = clock;
  assign buffer_3_reset = reset;
  assign buffer_3_auto_in_valid = cfar_auto_master_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_data = cfar_auto_master_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_last = cfar_auto_master_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_out_ready = widthAdapter_1_auto_in_ready; // @[LazyModule.scala 167:31]
  assign bus_clock = clock;
  assign bus_reset = reset;
  assign bus_auto_in_aw_valid = converter_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_id = converter_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_addr = converter_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_valid = converter_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_data = converter_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_strb = converter_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_last = converter_auto_out_w_bits_last; // @[LazyModule.scala 167:31]
  assign bus_auto_in_b_ready = converter_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_valid = converter_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_id = converter_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_addr = converter_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_size = converter_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_r_ready = converter_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_aw_ready = cfar_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_w_ready = cfar_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_b_valid = cfar_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_b_bits_id = cfar_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_ar_ready = cfar_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_r_valid = cfar_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_r_bits_id = cfar_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_2_r_bits_data = cfar_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_aw_ready = mag_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_w_ready = mag_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_b_valid = mag_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_b_bits_id = mag_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_ar_ready = mag_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_r_valid = mag_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_r_bits_id = mag_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_1_r_bits_data = mag_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_aw_ready = fft_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_w_ready = fft_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_b_valid = fft_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_b_bits_id = fft_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_ar_ready = fft_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_r_valid = fft_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_r_bits_id = fft_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_out_0_r_bits_data = fft_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign converter_auto_in_aw_valid = ioMem_0_aw_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_id = ioMem_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_addr = ioMem_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_valid = ioMem_0_w_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_data = ioMem_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_strb = ioMem_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_last = ioMem_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign converter_auto_in_b_ready = ioMem_0_b_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_valid = ioMem_0_ar_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_id = ioMem_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_addr = ioMem_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_size = ioMem_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_r_ready = ioMem_0_r_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_out_aw_ready = bus_auto_in_aw_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_w_ready = bus_auto_in_w_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_valid = bus_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_bits_resp = bus_auto_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_ar_ready = bus_auto_in_ar_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_valid = bus_auto_in_r_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_data = bus_auto_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_resp = bus_auto_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_last = bus_auto_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign converter_1_auto_in_valid = widthAdapter_1_auto_out_valid; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_data = widthAdapter_1_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_last = widthAdapter_1_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign converter_1_auto_out_ready = out_0_ready; // @[LazyModule.scala 167:31]
  assign converter_2_auto_in_valid = in_0_valid; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_data = in_0_bits_data; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_last = in_0_bits_last; // @[LazyModule.scala 167:57]
  assign converter_2_auto_out_ready = widthAdapter_auto_in_ready; // @[LazyModule.scala 167:31]
endmodule
module SRAM_depth_256_width_32_mem(
  input  [7:0]  R0_addr,
  input         R0_en,
  input         R0_clk,
  output [15:0] R0_data_real,
  output [15:0] R0_data_imag,
  input  [7:0]  W0_addr,
  input         W0_en,
  input         W0_clk,
  input  [15:0] W0_data_real,
  input  [15:0] W0_data_imag
);
  wire [7:0] SRAM_depth_256_width_32_mem_ext_R0_addr;
  wire  SRAM_depth_256_width_32_mem_ext_R0_en;
  wire  SRAM_depth_256_width_32_mem_ext_R0_clk;
  wire [31:0] SRAM_depth_256_width_32_mem_ext_R0_data;
  wire [7:0] SRAM_depth_256_width_32_mem_ext_W0_addr;
  wire  SRAM_depth_256_width_32_mem_ext_W0_en;
  wire  SRAM_depth_256_width_32_mem_ext_W0_clk;
  wire [31:0] SRAM_depth_256_width_32_mem_ext_W0_data;
  SRAM_depth_256_width_32_mem_ext SRAM_depth_256_width_32_mem_ext (
    .R0_addr(SRAM_depth_256_width_32_mem_ext_R0_addr),
    .R0_en(SRAM_depth_256_width_32_mem_ext_R0_en),
    .R0_clk(SRAM_depth_256_width_32_mem_ext_R0_clk),
    .R0_data(SRAM_depth_256_width_32_mem_ext_R0_data),
    .W0_addr(SRAM_depth_256_width_32_mem_ext_W0_addr),
    .W0_en(SRAM_depth_256_width_32_mem_ext_W0_en),
    .W0_clk(SRAM_depth_256_width_32_mem_ext_W0_clk),
    .W0_data(SRAM_depth_256_width_32_mem_ext_W0_data)
  );
  assign SRAM_depth_256_width_32_mem_ext_R0_clk = R0_clk;
  assign SRAM_depth_256_width_32_mem_ext_R0_en = R0_en;
  assign SRAM_depth_256_width_32_mem_ext_R0_addr = R0_addr;
  assign R0_data_imag = SRAM_depth_256_width_32_mem_ext_R0_data[15:0];
  assign R0_data_real = SRAM_depth_256_width_32_mem_ext_R0_data[31:16];
  assign SRAM_depth_256_width_32_mem_ext_W0_clk = W0_clk;
  assign SRAM_depth_256_width_32_mem_ext_W0_en = W0_en;
  assign SRAM_depth_256_width_32_mem_ext_W0_addr = W0_addr;
  assign SRAM_depth_256_width_32_mem_ext_W0_data = {W0_data_real,W0_data_imag};
endmodule
